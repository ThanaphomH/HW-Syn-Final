// *************************************************************
// Created by David J. Marion aka FPGA Dude
// A ROM containing patterns for ASCII values.
//
// Non-printable characters 00 - 1f, and 7f
// Printable characters 20 - 7e
//
// Not all character ROMs have been patterned.
// Only numbers, capital letters, some spec chars. 
//		Numbers       30 - 39
//   	Letters       41 - 5a 
//      (smiley face)   01
//		(space)         20
//		   .            2e
// 		   :            3a
//		   |	        7c	
//
// The 7-bit ASCII code for each character is used as
// the MSB of the address. The 4-bit LSB is the row value.
// *************************************************************

module thai_rom(
        input clk, 
        input wire [11:0] addr,
        output reg [7:0] data
    );

    (* rom_style = "block" *) 

    reg [10:0] addr_reg;
    
    always @(posedge clk)
        addr_reg <= addr;
        
    always @*
        case(addr_reg)
           // code x2D (-)
        12'h2D0: data = 8'b00000000;	//         
        12'h2D1: data = 8'b00000000;	//         
        12'h2D2: data = 8'b00000000;	//  
        12'h2D3: data = 8'b00000000;	// 
        12'h2D4: data = 8'b00000000;	// 
        12'h2D5: data = 8'b00000000;	// 
        12'h2D6: data = 8'b00000000;	// 
        12'h2D7: data = 8'b11111110;	// ******* 
        12'h2D8: data = 8'b11111110;	// ******* 
        12'h2D9: data = 8'b00000000;	// 
        12'h2Da: data = 8'b00000000;	//         
        12'h2Db: data = 8'b00000000;	//         
        12'h2Dc: data = 8'b00000000;	//         
        12'h2Dd: data = 8'b00000000;	//         
        12'h2De: data = 8'b00000000;	//         
        12'h2Df: data = 8'b00000000;	//  
             
    // code xe01 (ก)
        12'h010: data = 8'b00000000;	//         
        12'h011: data = 8'b00000000;	//         
        12'h012: data = 8'b00000000;	//         
        12'h013: data = 8'b00111100;	//   ****  
        12'h014: data = 8'b11000010;	// **    * 
        12'h015: data = 8'b11000010;	// **    * 
        12'h016: data = 8'b11000010;	// **    * 
        12'h017: data = 8'b11000010;	// **    * 
        12'h018: data = 8'b11000010;	// **    * 
        12'h019: data = 8'b11000010;	// **    * 
        12'h01a: data = 8'b00000000;	//         
        12'h01b: data = 8'b00000000;	//         
        12'h01c: data = 8'b00000000;	//         
        12'h01d: data = 8'b00000000;	//         
        12'h01e: data = 8'b00000000;	//         
        12'h01f: data = 8'b00000000;	//         

    // code xe02 (ข)
        12'h020: data = 8'b00000000;	//         
        12'h021: data = 8'b00000000;	//         
        12'h022: data = 8'b00000000;	//         
        12'h023: data = 8'b11001000;	// **  *   
        12'h024: data = 8'b11001000;	// **  *   
        12'h025: data = 8'b11001000;	// **  *   
        12'h026: data = 8'b11001000;	// **  *   
        12'h027: data = 8'b11001000;	// **  *   
        12'h028: data = 8'b11001000;	// **  *   
        12'h029: data = 8'b00110000;	//   **    
        12'h02a: data = 8'b00000000;	//         
        12'h02b: data = 8'b00000000;	//         
        12'h02c: data = 8'b00000000;	//         
        12'h02d: data = 8'b00000000;	//         
        12'h02e: data = 8'b00000000;	//         
        12'h02f: data = 8'b00000000;	//         

    // code xe03 (ฃ)
        12'h030: data = 8'b00000000;	//         
        12'h031: data = 8'b00000000;	//         
        12'h032: data = 8'b00000000;	//         
        12'h033: data = 8'b10000100;	// *    *  
        12'h034: data = 8'b00100100;	//   *  *  
        12'h035: data = 8'b00100100;	//   *  *  
        12'h036: data = 8'b00100100;	//   *  *  
        12'h037: data = 8'b00100100;	//   *  *  
        12'h038: data = 8'b00100100;	//   *  *  
        12'h039: data = 8'b00011000;	//    **   
        12'h03a: data = 8'b00000000;	//         
        12'h03b: data = 8'b00000000;	//         
        12'h03c: data = 8'b00000000;	//         
        12'h03d: data = 8'b00000000;	//         
        12'h03e: data = 8'b00000000;	//         
        12'h03f: data = 8'b00000000;	//         

    // code xe04 (ค)
        12'h040: data = 8'b00000000;	//         
        12'h041: data = 8'b00000000;	//         
        12'h042: data = 8'b00000000;	//         
        12'h043: data = 8'b00111100;	//   ****  
        12'h044: data = 8'b11000010;	// **    * 
        12'h045: data = 8'b11000010;	// **    * 
        12'h046: data = 8'b11000010;	// **    * 
        12'h047: data = 8'b11110010;	// ****  * 
        12'h048: data = 8'b11000010;	// **    * 
        12'h049: data = 8'b11000010;	// **    * 
        12'h04a: data = 8'b00000000;	//         
        12'h04b: data = 8'b00000000;	//         
        12'h04c: data = 8'b00000000;	//         
        12'h04d: data = 8'b00000000;	//         
        12'h04e: data = 8'b00000000;	//         
        12'h04f: data = 8'b00000000;	//         

    // code xe05 (ฅ)
        12'h050: data = 8'b00000000;	//         
        12'h051: data = 8'b00000000;	//         
        12'h052: data = 8'b00000000;	//         
        12'h053: data = 8'b00100100;	//   *  *  
        12'h054: data = 8'b11000010;	// **    * 
        12'h055: data = 8'b11000010;	// **    * 
        12'h056: data = 8'b11000010;	// **    * 
        12'h057: data = 8'b11110010;	// ****  * 
        12'h058: data = 8'b11000010;	// **    * 
        12'h059: data = 8'b11000010;	// **    * 
        12'h05a: data = 8'b00000000;	//         
        12'h05b: data = 8'b00000000;	//         
        12'h05c: data = 8'b00000000;	//         
        12'h05d: data = 8'b00000000;	//         
        12'h05e: data = 8'b00000000;	//         
        12'h05f: data = 8'b00000000;	//         

    // code xe06 (ฆ)
        12'h060: data = 8'b00000000;	//         
        12'h061: data = 8'b00000000;	//         
        12'h062: data = 8'b00000000;	//         
        12'h063: data = 8'b10000010;	// *     * 
        12'h064: data = 8'b00100010;	//   *   * 
        12'h065: data = 8'b00100010;	//   *   * 
        12'h066: data = 8'b00100010;	//   *   * 
        12'h067: data = 8'b00100010;	//   *   * 
        12'h068: data = 8'b01110000;	//  ***    
        12'h069: data = 8'b00100100;	//   *  *  
        12'h06a: data = 8'b00000000;	//         
        12'h06b: data = 8'b00000000;	//         
        12'h06c: data = 8'b00000000;	//         
        12'h06d: data = 8'b00000000;	//         
        12'h06e: data = 8'b00000000;	//         
        12'h06f: data = 8'b00000000;	//         

    // code xe07 (ง)
        12'h070: data = 8'b00000000;	//         
        12'h071: data = 8'b00000000;	//         
        12'h072: data = 8'b00000000;	//         
        12'h073: data = 8'b00011000;	//    **   
        12'h074: data = 8'b00001000;	//     *   
        12'h075: data = 8'b00001000;	//     *   
        12'h076: data = 8'b11001000;	// **  *   
        12'h077: data = 8'b11001000;	// **  *   
        12'h078: data = 8'b11001000;	// **  *   
        12'h079: data = 8'b00110000;	//   **    
        12'h07a: data = 8'b00000000;	//         
        12'h07b: data = 8'b00000000;	//         
        12'h07c: data = 8'b00000000;	//         
        12'h07d: data = 8'b00000000;	//         
        12'h07e: data = 8'b00000000;	//         
        12'h07f: data = 8'b00000000;	//         

    // code xe08 (จ)
        12'h080: data = 8'b00000000;	//         
        12'h081: data = 8'b00000000;	//         
        12'h082: data = 8'b00000000;	//         
        12'h083: data = 8'b00111100;	//   ****  
        12'h084: data = 8'b00000010;	//       * 
        12'h085: data = 8'b11000010;	// **    * 
        12'h086: data = 8'b00000010;	//       * 
        12'h087: data = 8'b00001110;	//     *** 
        12'h088: data = 8'b00000010;	//       * 
        12'h089: data = 8'b00000010;	//       * 
        12'h08a: data = 8'b00000000;	//         
        12'h08b: data = 8'b00000000;	//         
        12'h08c: data = 8'b00000000;	//         
        12'h08d: data = 8'b00000000;	//         
        12'h08e: data = 8'b00000000;	//         
        12'h08f: data = 8'b00000000;	//         

    // code xe09 (ฉ)
        12'h090: data = 8'b00000000;	//         
        12'h091: data = 8'b00000000;	//         
        12'h092: data = 8'b00000000;	//         
        12'h093: data = 8'b00111100;	//   ****  
        12'h094: data = 8'b11000000;	// **      
        12'h095: data = 8'b11000010;	// **    * 
        12'h096: data = 8'b00000010;	//       * 
        12'h097: data = 8'b11000010;	// **    * 
        12'h098: data = 8'b11001111;	// **  ****
        12'h099: data = 8'b00100010;	//   *   * 
        12'h09a: data = 8'b00000000;	//         
        12'h09b: data = 8'b00000000;	//         
        12'h09c: data = 8'b00000000;	//         
        12'h09d: data = 8'b00000000;	//         
        12'h09e: data = 8'b00000000;	//         
        12'h09f: data = 8'b00000000;	//         

    // code xe0a (ช)
        12'h0a0: data = 8'b00000000;	//         
        12'h0a1: data = 8'b00000000;	//         
        12'h0a2: data = 8'b00000000;	//         
        12'h0a3: data = 8'b11001000;	// **  *   
        12'h0a4: data = 8'b11110000;	// ****    
        12'h0a5: data = 8'b11000000;	// **      
        12'h0a6: data = 8'b11001000;	// **  *   
        12'h0a7: data = 8'b11001000;	// **  *   
        12'h0a8: data = 8'b01001000;	//  *  *   
        12'h0a9: data = 8'b00110000;	//   **    
        12'h0aa: data = 8'b00000000;	//         
        12'h0ab: data = 8'b00000000;	//         
        12'h0ac: data = 8'b00000000;	//         
        12'h0ad: data = 8'b00000000;	//         
        12'h0ae: data = 8'b00000000;	//         
        12'h0af: data = 8'b00000000;	//         

    // code xe0b (ซ)
        12'h0b0: data = 8'b00000000;	//         
        12'h0b1: data = 8'b00000000;	//         
        12'h0b2: data = 8'b00000000;	//         
        12'h0b3: data = 8'b10000100;	// *    *  
        12'h0b4: data = 8'b00011000;	//    **   
        12'h0b5: data = 8'b00111000;	//   ***   
        12'h0b6: data = 8'b00100100;	//   *  *  
        12'h0b7: data = 8'b00100100;	//   *  *  
        12'h0b8: data = 8'b00100100;	//   *  *  
        12'h0b9: data = 8'b00011000;	//    **   
        12'h0ba: data = 8'b00000000;	//         
        12'h0bb: data = 8'b00000000;	//         
        12'h0bc: data = 8'b00000000;	//         
        12'h0bd: data = 8'b00000000;	//         
        12'h0be: data = 8'b00000000;	//         
        12'h0bf: data = 8'b00000000;	//         

    // code xe0c (ฌ)
        12'h0c0: data = 8'b00000000;	//         
        12'h0c1: data = 8'b00000000;	//         
        12'h0c2: data = 8'b00000000;	//         
        12'h0c3: data = 8'b00111100;	//   ****  
        12'h0c4: data = 8'b11000010;	// **    * 
        12'h0c5: data = 8'b11000010;	// **    * 
        12'h0c6: data = 8'b11000010;	// **    * 
        12'h0c7: data = 8'b11000010;	// **    * 
        12'h0c8: data = 8'b11000111;	// **   ***
        12'h0c9: data = 8'b11100010;	// ***   * 
        12'h0ca: data = 8'b00000000;	//         
        12'h0cb: data = 8'b00000000;	//         
        12'h0cc: data = 8'b00000000;	//         
        12'h0cd: data = 8'b00000000;	//         
        12'h0ce: data = 8'b00000000;	//         
        12'h0cf: data = 8'b00000000;	//         

    // code xe0d (ญ)
        12'h0d0: data = 8'b00000000;	//         
        12'h0d1: data = 8'b00000000;	//         
        12'h0d2: data = 8'b00000000;	//         
        12'h0d3: data = 8'b00111100;	//   ****  
        12'h0d4: data = 8'b11000010;	// **    * 
        12'h0d5: data = 8'b11000010;	// **    * 
        12'h0d6: data = 8'b11000010;	// **    * 
        12'h0d7: data = 8'b11000010;	// **    * 
        12'h0d8: data = 8'b11000001;	// **     *
        12'h0d9: data = 8'b11100000;	// ***     
        12'h0da: data = 8'b00000001;	//        *
        12'h0db: data = 8'b00000000;	//         
        12'h0dc: data = 8'b00000000;	//         
        12'h0dd: data = 8'b00000000;	//         
        12'h0de: data = 8'b00000000;	//         
        12'h0df: data = 8'b00000000;	//         

    // code xe0e (ฎ)
        12'h0e0: data = 8'b00000000;	//         
        12'h0e1: data = 8'b00000000;	//         
        12'h0e2: data = 8'b00000000;	//         
        12'h0e3: data = 8'b00111100;	//   ****  
        12'h0e4: data = 8'b11000010;	// **    * 
        12'h0e5: data = 8'b11000010;	// **    * 
        12'h0e6: data = 8'b11000010;	// **    * 
        12'h0e7: data = 8'b11000010;	// **    * 
        12'h0e8: data = 8'b11000010;	// **    * 
        12'h0e9: data = 8'b11000010;	// **    * 
        12'h0ea: data = 8'b00000010;	//       * 
        12'h0eb: data = 8'b00100100;	//   *  *  
        12'h0ec: data = 8'b00000000;	//         
        12'h0ed: data = 8'b00000000;	//         
        12'h0ee: data = 8'b00000000;	//         
        12'h0ef: data = 8'b00000000;	//         

    // code xe0f (ฏ)
        12'h0f0: data = 8'b00000000;	//         
        12'h0f1: data = 8'b00000000;	//         
        12'h0f2: data = 8'b00000000;	//         
        12'h0f3: data = 8'b00111100;	//   ****  
        12'h0f4: data = 8'b11000010;	// **    * 
        12'h0f5: data = 8'b11000010;	// **    * 
        12'h0f6: data = 8'b11000010;	// **    * 
        12'h0f7: data = 8'b11000010;	// **    * 
        12'h0f8: data = 8'b11000010;	// **    * 
        12'h0f9: data = 8'b11000010;	// **    * 
        12'h0fa: data = 8'b00000110;	//      ** 
        12'h0fb: data = 8'b00000010;	//       * 
        12'h0fc: data = 8'b00000000;	//         
        12'h0fd: data = 8'b00000000;	//         
        12'h0fe: data = 8'b00000000;	//         
        12'h0ff: data = 8'b00000000;	//         

    // code xe10 (ฐ)
        12'h100: data = 8'b00000000;	//         
        12'h101: data = 8'b00000000;	//         
        12'h102: data = 8'b00000000;	//         
        12'h103: data = 8'b00111110;	//   ***** 
        12'h104: data = 8'b00000010;	//       * 
        12'h105: data = 8'b00000010;	//       * 
        12'h106: data = 8'b00000010;	//       * 
        12'h107: data = 8'b00001110;	//     *** 
        12'h108: data = 8'b00000010;	//       * 
        12'h109: data = 8'b00000010;	//       * 
        12'h10a: data = 8'b00000000;	//         
        12'h10b: data = 8'b00000000;	//         
        12'h10c: data = 8'b00000000;	//         
        12'h10d: data = 8'b00000000;	//         
        12'h10e: data = 8'b00000000;	//         
        12'h10f: data = 8'b00000000;	//         

    // code xe11 (ฑ)
        12'h110: data = 8'b00000000;	//         
        12'h111: data = 8'b00000000;	//         
        12'h112: data = 8'b00000000;	//         
        12'h113: data = 8'b10000010;	// *     * 
        12'h114: data = 8'b00100001;	//   *    *
        12'h115: data = 8'b00100001;	//   *    *
        12'h116: data = 8'b00110001;	//   **   *
        12'h117: data = 8'b00100001;	//   *    *
        12'h118: data = 8'b00100001;	//   *    *
        12'h119: data = 8'b00100001;	//   *    *
        12'h11a: data = 8'b00000000;	//         
        12'h11b: data = 8'b00000000;	//         
        12'h11c: data = 8'b00000000;	//         
        12'h11d: data = 8'b00000000;	//         
        12'h11e: data = 8'b00000000;	//         
        12'h11f: data = 8'b00000000;	//         

    // code xe12 (ฒ)
        12'h120: data = 8'b00000000;	//         
        12'h121: data = 8'b00000000;	//         
        12'h122: data = 8'b00000000;	//         
        12'h123: data = 8'b00100100;	//   *  *  
        12'h124: data = 8'b11000010;	// **    * 
        12'h125: data = 8'b11000010;	// **    * 
        12'h126: data = 8'b11000010;	// **    * 
        12'h127: data = 8'b11000010;	// **    * 
        12'h128: data = 8'b11000111;	// **   ***
        12'h129: data = 8'b00100010;	//   *   * 
        12'h12a: data = 8'b00000000;	//         
        12'h12b: data = 8'b00000000;	//         
        12'h12c: data = 8'b00000000;	//         
        12'h12d: data = 8'b00000000;	//         
        12'h12e: data = 8'b00000000;	//         
        12'h12f: data = 8'b00000000;	//         

    // code xe13 (ณ)
        12'h130: data = 8'b00000000;	//         
        12'h131: data = 8'b00000000;	//         
        12'h132: data = 8'b00000000;	//         
        12'h133: data = 8'b00111100;	//   ****  
        12'h134: data = 8'b11000010;	// **    * 
        12'h135: data = 8'b11000010;	// **    * 
        12'h136: data = 8'b11000010;	// **    * 
        12'h137: data = 8'b11000010;	// **    * 
        12'h138: data = 8'b11000010;	// **    * 
        12'h139: data = 8'b11100001;	// ***    *
        12'h13a: data = 8'b00000000;	//         
        12'h13b: data = 8'b00000000;	//         
        12'h13c: data = 8'b00000000;	//         
        12'h13d: data = 8'b00000000;	//         
        12'h13e: data = 8'b00000000;	//         
        12'h13f: data = 8'b00000000;	//         

    // code xe14 (ด)
        12'h140: data = 8'b00000000;	//         
        12'h141: data = 8'b00000000;	//         
        12'h142: data = 8'b00000000;	//         
        12'h143: data = 8'b00111100;	//   ****  
        12'h144: data = 8'b11000010;	// **    * 
        12'h145: data = 8'b11000010;	// **    * 
        12'h146: data = 8'b11000010;	// **    * 
        12'h147: data = 8'b11000010;	// **    * 
        12'h148: data = 8'b11000010;	// **    * 
        12'h149: data = 8'b00110010;	//   **  * 
        12'h14a: data = 8'b00000000;	//         
        12'h14b: data = 8'b00000000;	//         
        12'h14c: data = 8'b00000000;	//         
        12'h14d: data = 8'b00000000;	//         
        12'h14e: data = 8'b00000000;	//         
        12'h14f: data = 8'b00000000;	//         

    // code xe15 (ต)
        12'h150: data = 8'b00000000;	//         
        12'h151: data = 8'b00000000;	//         
        12'h152: data = 8'b00000000;	//         
        12'h153: data = 8'b00100100;	//   *  *  
        12'h154: data = 8'b11000010;	// **    * 
        12'h155: data = 8'b11000010;	// **    * 
        12'h156: data = 8'b11000010;	// **    * 
        12'h157: data = 8'b11000010;	// **    * 
        12'h158: data = 8'b11000010;	// **    * 
        12'h159: data = 8'b00110010;	//   **  * 
        12'h15a: data = 8'b00000000;	//         
        12'h15b: data = 8'b00000000;	//         
        12'h15c: data = 8'b00000000;	//         
        12'h15d: data = 8'b00000000;	//         
        12'h15e: data = 8'b00000000;	//         
        12'h15f: data = 8'b00000000;	//         

    // code xe16 (ถ)
        12'h160: data = 8'b00000000;	//         
        12'h161: data = 8'b00000000;	//         
        12'h162: data = 8'b00000000;	//         
        12'h163: data = 8'b00111100;	//   ****  
        12'h164: data = 8'b11000010;	// **    * 
        12'h165: data = 8'b11000010;	// **    * 
        12'h166: data = 8'b11000010;	// **    * 
        12'h167: data = 8'b11000010;	// **    * 
        12'h168: data = 8'b11000010;	// **    * 
        12'h169: data = 8'b11100010;	// ***   * 
        12'h16a: data = 8'b00000000;	//         
        12'h16b: data = 8'b00000000;	//         
        12'h16c: data = 8'b00000000;	//         
        12'h16d: data = 8'b00000000;	//         
        12'h16e: data = 8'b00000000;	//         
        12'h16f: data = 8'b00000000;	//         

    // code xe17 (ท)
        12'h170: data = 8'b00000000;	//         
        12'h171: data = 8'b00000000;	//         
        12'h172: data = 8'b00000000;	//         
        12'h173: data = 8'b11000100;	// **   *  
        12'h174: data = 8'b11000010;	// **    * 
        12'h175: data = 8'b11100010;	// ***   * 
        12'h176: data = 8'b11000010;	// **    * 
        12'h177: data = 8'b11000010;	// **    * 
        12'h178: data = 8'b11000010;	// **    * 
        12'h179: data = 8'b11000010;	// **    * 
        12'h17a: data = 8'b00000000;	//         
        12'h17b: data = 8'b00000000;	//         
        12'h17c: data = 8'b00000000;	//         
        12'h17d: data = 8'b00000000;	//         
        12'h17e: data = 8'b00000000;	//         
        12'h17f: data = 8'b00000000;	//         

    // code xe18 (ธ)
        12'h180: data = 8'b00000000;	//         
        12'h181: data = 8'b00000000;	//         
        12'h182: data = 8'b00000000;	//         
        12'h183: data = 8'b00111110;	//   ***** 
        12'h184: data = 8'b11000000;	// **      
        12'h185: data = 8'b00000000;	//         
        12'h186: data = 8'b00111100;	//   ****  
        12'h187: data = 8'b00000010;	//       * 
        12'h188: data = 8'b11000010;	// **    * 
        12'h189: data = 8'b11111100;	// ******  
        12'h18a: data = 8'b00000000;	//         
        12'h18b: data = 8'b00000000;	//         
        12'h18c: data = 8'b00000000;	//         
        12'h18d: data = 8'b00000000;	//         
        12'h18e: data = 8'b00000000;	//         
        12'h18f: data = 8'b00000000;	//         

    // code xe19 (น)
        12'h190: data = 8'b00000000;	//         
        12'h191: data = 8'b00000000;	//         
        12'h192: data = 8'b00000000;	//         
        12'h193: data = 8'b11000010;	// **    * 
        12'h194: data = 8'b11000010;	// **    * 
        12'h195: data = 8'b11000010;	// **    * 
        12'h196: data = 8'b11000010;	// **    * 
        12'h197: data = 8'b11000010;	// **    * 
        12'h198: data = 8'b01000011;	//  *    **
        12'h199: data = 8'b00100010;	//   *   * 
        12'h19a: data = 8'b00000000;	//         
        12'h19b: data = 8'b00000000;	//         
        12'h19c: data = 8'b00000000;	//         
        12'h19d: data = 8'b00000000;	//         
        12'h19e: data = 8'b00000000;	//         
        12'h19f: data = 8'b00000000;	//         

    // code xe1a (บ)
        12'h1a0: data = 8'b00000000;	//         
        12'h1a1: data = 8'b00000000;	//         
        12'h1a2: data = 8'b00000000;	//         
        12'h1a3: data = 8'b11000010;	// **    * 
        12'h1a4: data = 8'b11000010;	// **    * 
        12'h1a5: data = 8'b11000010;	// **    * 
        12'h1a6: data = 8'b11000010;	// **    * 
        12'h1a7: data = 8'b11000010;	// **    * 
        12'h1a8: data = 8'b11000010;	// **    * 
        12'h1a9: data = 8'b00111100;	//   ****  
        12'h1aa: data = 8'b00000000;	//         
        12'h1ab: data = 8'b00000000;	//         
        12'h1ac: data = 8'b00000000;	//         
        12'h1ad: data = 8'b00000000;	//         
        12'h1ae: data = 8'b00000000;	//         
        12'h1af: data = 8'b00000000;	//         

    // code xe1b (ป)
        12'h1b0: data = 8'b00000000;	//         
        12'h1b1: data = 8'b00000010;	//       * 
        12'h1b2: data = 8'b00000010;	//       * 
        12'h1b3: data = 8'b00000010;	//       * 
        12'h1b4: data = 8'b11000010;	// **    * 
        12'h1b5: data = 8'b11000010;	// **    * 
        12'h1b6: data = 8'b11000010;	// **    * 
        12'h1b7: data = 8'b11000010;	// **    * 
        12'h1b8: data = 8'b11000010;	// **    * 
        12'h1b9: data = 8'b00111100;	//   ****  
        12'h1ba: data = 8'b00000000;	//         
        12'h1bb: data = 8'b00000000;	//         
        12'h1bc: data = 8'b00000000;	//         
        12'h1bd: data = 8'b00000000;	//         
        12'h1be: data = 8'b00000000;	//         
        12'h1bf: data = 8'b00000000;	//         

    // code xe1c (ผ)
        12'h1c0: data = 8'b00000000;	//         
        12'h1c1: data = 8'b00000000;	//         
        12'h1c2: data = 8'b00000000;	//         
        12'h1c3: data = 8'b00100010;	//   *   * 
        12'h1c4: data = 8'b11000010;	// **    * 
        12'h1c5: data = 8'b11000010;	// **    * 
        12'h1c6: data = 8'b11000010;	// **    * 
        12'h1c7: data = 8'b11000010;	// **    * 
        12'h1c8: data = 8'b11000010;	// **    * 
        12'h1c9: data = 8'b00100100;	//   *  *  
        12'h1ca: data = 8'b00000000;	//         
        12'h1cb: data = 8'b00000000;	//         
        12'h1cc: data = 8'b00000000;	//         
        12'h1cd: data = 8'b00000000;	//         
        12'h1ce: data = 8'b00000000;	//         
        12'h1cf: data = 8'b00000000;	//         

    // code xe1d (ฝ)
        12'h1d0: data = 8'b00000000;	//         
        12'h1d1: data = 8'b00000010;	//       * 
        12'h1d2: data = 8'b00000010;	//       * 
        12'h1d3: data = 8'b00100010;	//   *   * 
        12'h1d4: data = 8'b11000010;	// **    * 
        12'h1d5: data = 8'b11000010;	// **    * 
        12'h1d6: data = 8'b11000010;	// **    * 
        12'h1d7: data = 8'b11000010;	// **    * 
        12'h1d8: data = 8'b11000010;	// **    * 
        12'h1d9: data = 8'b00100100;	//   *  *  
        12'h1da: data = 8'b00000000;	//         
        12'h1db: data = 8'b00000000;	//         
        12'h1dc: data = 8'b00000000;	//         
        12'h1dd: data = 8'b00000000;	//         
        12'h1de: data = 8'b00000000;	//         
        12'h1df: data = 8'b00000000;	//         

    // code xe1e (พ)
        12'h1e0: data = 8'b00000000;	//         
        12'h1e1: data = 8'b00000000;	//         
        12'h1e2: data = 8'b00000000;	//         
        12'h1e3: data = 8'b11000010;	// **    * 
        12'h1e4: data = 8'b11000010;	// **    * 
        12'h1e5: data = 8'b11000010;	// **    * 
        12'h1e6: data = 8'b11000010;	// **    * 
        12'h1e7: data = 8'b11000010;	// **    * 
        12'h1e8: data = 8'b11000010;	// **    * 
        12'h1e9: data = 8'b00100100;	//   *  *  
        12'h1ea: data = 8'b00000000;	//         
        12'h1eb: data = 8'b00000000;	//         
        12'h1ec: data = 8'b00000000;	//         
        12'h1ed: data = 8'b00000000;	//         
        12'h1ee: data = 8'b00000000;	//         
        12'h1ef: data = 8'b00000000;	//         

    // code xe1f (ฟ)
        12'h1f0: data = 8'b00000000;	//         
        12'h1f1: data = 8'b00000010;	//       * 
        12'h1f2: data = 8'b00000010;	//       * 
        12'h1f3: data = 8'b00000010;	//       * 
        12'h1f4: data = 8'b11000010;	// **    * 
        12'h1f5: data = 8'b11000010;	// **    * 
        12'h1f6: data = 8'b11000010;	// **    * 
        12'h1f7: data = 8'b11000010;	// **    * 
        12'h1f8: data = 8'b11000010;	// **    * 
        12'h1f9: data = 8'b00100100;	//   *  *  
        12'h1fa: data = 8'b00000000;	//         
        12'h1fb: data = 8'b00000000;	//         
        12'h1fc: data = 8'b00000000;	//         
        12'h1fd: data = 8'b00000000;	//         
        12'h1fe: data = 8'b00000000;	//         
        12'h1ff: data = 8'b00000000;	//         

    // code xe20 (ภ)
        12'h200: data = 8'b00000000;	//         
        12'h201: data = 8'b00000000;	//         
        12'h202: data = 8'b00000000;	//         
        12'h203: data = 8'b00011110;	//    **** 
        12'h204: data = 8'b00100001;	//   *    *
        12'h205: data = 8'b00100001;	//   *    *
        12'h206: data = 8'b00100001;	//   *    *
        12'h207: data = 8'b00100001;	//   *    *
        12'h208: data = 8'b00100001;	//   *    *
        12'h209: data = 8'b11100001;	// ***    *
        12'h20a: data = 8'b00000000;	//         
        12'h20b: data = 8'b00000000;	//         
        12'h20c: data = 8'b00000000;	//         
        12'h20d: data = 8'b00000000;	//         
        12'h20e: data = 8'b00000000;	//         
        12'h20f: data = 8'b00000000;	//         

    // code xe21 (ม)
        12'h210: data = 8'b00000000;	//         
        12'h211: data = 8'b00000000;	//         
        12'h212: data = 8'b00000000;	//         
        12'h213: data = 8'b11100001;	// ***    *
        12'h214: data = 8'b00100001;	//   *    *
        12'h215: data = 8'b00100001;	//   *    *
        12'h216: data = 8'b00100001;	//   *    *
        12'h217: data = 8'b00100001;	//   *    *
        12'h218: data = 8'b11111001;	// *****  *
        12'h219: data = 8'b00100010;	//   *   * 
        12'h21a: data = 8'b00000000;	//         
        12'h21b: data = 8'b00000000;	//         
        12'h21c: data = 8'b00000000;	//         
        12'h21d: data = 8'b00000000;	//         
        12'h21e: data = 8'b00000000;	//         
        12'h21f: data = 8'b00000000;	//         

    // code xe22 (ย)
        12'h220: data = 8'b00000000;	//         
        12'h221: data = 8'b00000000;	//         
        12'h222: data = 8'b00000000;	//         
        12'h223: data = 8'b00100010;	//   *   * 
        12'h224: data = 8'b11000010;	// **    * 
        12'h225: data = 8'b00000010;	//       * 
        12'h226: data = 8'b00110010;	//   **  * 
        12'h227: data = 8'b11000010;	// **    * 
        12'h228: data = 8'b11000010;	// **    * 
        12'h229: data = 8'b00111100;	//   ****  
        12'h22a: data = 8'b00000000;	//         
        12'h22b: data = 8'b00000000;	//         
        12'h22c: data = 8'b00000000;	//         
        12'h22d: data = 8'b00000000;	//         
        12'h22e: data = 8'b00000000;	//         
        12'h22f: data = 8'b00000000;	//         

    // code xe23 (ร)
        12'h230: data = 8'b00000000;	//         
        12'h231: data = 8'b00000000;	//         
        12'h232: data = 8'b00000000;	//         
        12'h233: data = 8'b00111100;	//   ****  
        12'h234: data = 8'b11000000;	// **      
        12'h235: data = 8'b00000000;	//         
        12'h236: data = 8'b00111000;	//   ***   
        12'h237: data = 8'b00000100;	//      *  
        12'h238: data = 8'b00000100;	//      *  
        12'h239: data = 8'b00011000;	//    **   
        12'h23a: data = 8'b00000000;	//         
        12'h23b: data = 8'b00000000;	//         
        12'h23c: data = 8'b00000000;	//         
        12'h23d: data = 8'b00000000;	//         
        12'h23e: data = 8'b00000000;	//         
        12'h23f: data = 8'b00000000;	//         

    // code xe24 (ฤ)
        12'h240: data = 8'b00000000;	//         
        12'h241: data = 8'b00000000;	//         
        12'h242: data = 8'b00000000;	//         
        12'h243: data = 8'b00111100;	//   ****  
        12'h244: data = 8'b11000010;	// **    * 
        12'h245: data = 8'b11000010;	// **    * 
        12'h246: data = 8'b11000010;	// **    * 
        12'h247: data = 8'b11000010;	// **    * 
        12'h248: data = 8'b11000010;	// **    * 
        12'h249: data = 8'b11100010;	// ***   * 
        12'h24a: data = 8'b00000010;	//       * 
        12'h24b: data = 8'b00000010;	//       * 
        12'h24c: data = 8'b00000000;	//         
        12'h24d: data = 8'b00000000;	//         
        12'h24e: data = 8'b00000000;	//         
        12'h24f: data = 8'b00000000;	//         

    // code xe25 (ล)
        12'h250: data = 8'b00000000;	//         
        12'h251: data = 8'b00000000;	//         
        12'h252: data = 8'b00000000;	//         
        12'h253: data = 8'b11111100;	// ******  
        12'h254: data = 8'b00000010;	//       * 
        12'h255: data = 8'b00000010;	//       * 
        12'h256: data = 8'b00111110;	//   ***** 
        12'h257: data = 8'b11000010;	// **    * 
        12'h258: data = 8'b01000010;	//  *    * 
        12'h259: data = 8'b00100010;	//   *   * 
        12'h25a: data = 8'b00000000;	//         
        12'h25b: data = 8'b00000000;	//         
        12'h25c: data = 8'b00000000;	//         
        12'h25d: data = 8'b00000000;	//         
        12'h25e: data = 8'b00000000;	//         
        12'h25f: data = 8'b00000000;	//         

    // code xe26 (ฦ)
        12'h260: data = 8'b00000000;	//         
        12'h261: data = 8'b00000000;	//         
        12'h262: data = 8'b00000000;	//         
        12'h263: data = 8'b00011110;	//    **** 
        12'h264: data = 8'b00100001;	//   *    *
        12'h265: data = 8'b00100001;	//   *    *
        12'h266: data = 8'b00100001;	//   *    *
        12'h267: data = 8'b00100001;	//   *    *
        12'h268: data = 8'b00100001;	//   *    *
        12'h269: data = 8'b11100001;	// ***    *
        12'h26a: data = 8'b00000001;	//        *
        12'h26b: data = 8'b00000001;	//        *
        12'h26c: data = 8'b00000000;	//         
        12'h26d: data = 8'b00000000;	//         
        12'h26e: data = 8'b00000000;	//         
        12'h26f: data = 8'b00000000;	//         

    // code xe27 (ว)
        12'h270: data = 8'b00000000;	//         
        12'h271: data = 8'b00000000;	//         
        12'h272: data = 8'b00000000;	//         
        12'h273: data = 8'b11111000;	// *****   
        12'h274: data = 8'b00000100;	//      *  
        12'h275: data = 8'b00000100;	//      *  
        12'h276: data = 8'b00000100;	//      *  
        12'h277: data = 8'b00000100;	//      *  
        12'h278: data = 8'b00000100;	//      *  
        12'h279: data = 8'b00011000;	//    **   
        12'h27a: data = 8'b00000000;	//         
        12'h27b: data = 8'b00000000;	//         
        12'h27c: data = 8'b00000000;	//         
        12'h27d: data = 8'b00000000;	//         
        12'h27e: data = 8'b00000000;	//         
        12'h27f: data = 8'b00000000;	//         

    // code xe28 (ศ)
        12'h280: data = 8'b00000000;	//         
        12'h281: data = 8'b00000000;	//         
        12'h282: data = 8'b00000010;	//       * 
        12'h283: data = 8'b00111110;	//   ***** 
        12'h284: data = 8'b11000010;	// **    * 
        12'h285: data = 8'b11000010;	// **    * 
        12'h286: data = 8'b11000010;	// **    * 
        12'h287: data = 8'b11110010;	// ****  * 
        12'h288: data = 8'b11000010;	// **    * 
        12'h289: data = 8'b11000010;	// **    * 
        12'h28a: data = 8'b00000000;	//         
        12'h28b: data = 8'b00000000;	//         
        12'h28c: data = 8'b00000000;	//         
        12'h28d: data = 8'b00000000;	//         
        12'h28e: data = 8'b00000000;	//         
        12'h28f: data = 8'b00000000;	//         

    // code xe29 (ษ)
        12'h290: data = 8'b00000000;	//         
        12'h291: data = 8'b00000000;	//         
        12'h292: data = 8'b00000000;	//         
        12'h293: data = 8'b11000010;	// **    * 
        12'h294: data = 8'b11000010;	// **    * 
        12'h295: data = 8'b11000010;	// **    * 
        12'h296: data = 8'b11001110;	// **  *** 
        12'h297: data = 8'b11000010;	// **    * 
        12'h298: data = 8'b11000010;	// **    * 
        12'h299: data = 8'b00111100;	//   ****  
        12'h29a: data = 8'b00000000;	//         
        12'h29b: data = 8'b00000000;	//         
        12'h29c: data = 8'b00000000;	//         
        12'h29d: data = 8'b00000000;	//         
        12'h29e: data = 8'b00000000;	//         
        12'h29f: data = 8'b00000000;	//         

    // code xe2a (ส)
        12'h2a0: data = 8'b00000000;	//         
        12'h2a1: data = 8'b00000000;	//         
        12'h2a2: data = 8'b00000010;	//       * 
        12'h2a3: data = 8'b11111110;	// ******* 
        12'h2a4: data = 8'b00000010;	//       * 
        12'h2a5: data = 8'b00000010;	//       * 
        12'h2a6: data = 8'b00111110;	//   ***** 
        12'h2a7: data = 8'b11000010;	// **    * 
        12'h2a8: data = 8'b01000010;	//  *    * 
        12'h2a9: data = 8'b00100010;	//   *   * 
        12'h2aa: data = 8'b00000000;	//         
        12'h2ab: data = 8'b00000000;	//         
        12'h2ac: data = 8'b00000000;	//         
        12'h2ad: data = 8'b00000000;	//         
        12'h2ae: data = 8'b00000000;	//         
        12'h2af: data = 8'b00000000;	//         

    // code xe2b (ห)
        12'h2b0: data = 8'b00000000;	//         
        12'h2b1: data = 8'b00000000;	//         
        12'h2b2: data = 8'b00000000;	//         
        12'h2b3: data = 8'b00000000;	//         
        12'h2b4: data = 8'b11000010;	// **    * 
        12'h2b5: data = 8'b11000010;	// **    * 
        12'h2b6: data = 8'b11000100;	// **   *  
        12'h2b7: data = 8'b11000010;	// **    * 
        12'h2b8: data = 8'b11100010;	// ***   * 
        12'h2b9: data = 8'b11000010;	// **    * 
        12'h2ba: data = 8'b00000000;	//         
        12'h2bb: data = 8'b00000000;	//         
        12'h2bc: data = 8'b00000000;	//         
        12'h2bd: data = 8'b00000000;	//         
        12'h2be: data = 8'b00000000;	//         
        12'h2bf: data = 8'b00000000;	//         

    // code xe2c (ฬ)
        12'h2c0: data = 8'b00000000;	//         
        12'h2c1: data = 8'b00000000;	//         
        12'h2c2: data = 8'b00000000;	//         
        12'h2c3: data = 8'b11000010;	// **    * 
        12'h2c4: data = 8'b11000100;	// **   *  
        12'h2c5: data = 8'b11000100;	// **   *  
        12'h2c6: data = 8'b11000010;	// **    * 
        12'h2c7: data = 8'b11000010;	// **    * 
        12'h2c8: data = 8'b01000010;	//  *    * 
        12'h2c9: data = 8'b00100100;	//   *  *  
        12'h2ca: data = 8'b00000000;	//         
        12'h2cb: data = 8'b00000000;	//         
        12'h2cc: data = 8'b00000000;	//         
        12'h2cd: data = 8'b00000000;	//         
        12'h2ce: data = 8'b00000000;	//         
        12'h2cf: data = 8'b00000000;	//         

    // code xe2d (อ)
        12'h2d0: data = 8'b00000000;	//         
        12'h2d1: data = 8'b00000000;	//         
        12'h2d2: data = 8'b00000000;	//         
        12'h2d3: data = 8'b11111100;	// ******  
        12'h2d4: data = 8'b00000010;	//       * 
        12'h2d5: data = 8'b00000010;	//       * 
        12'h2d6: data = 8'b11100010;	// ***   * 
        12'h2d7: data = 8'b11000010;	// **    * 
        12'h2d8: data = 8'b11000010;	// **    * 
        12'h2d9: data = 8'b00111100;	//   ****  
        12'h2da: data = 8'b00000000;	//         
        12'h2db: data = 8'b00000000;	//         
        12'h2dc: data = 8'b00000000;	//         
        12'h2dd: data = 8'b00000000;	//         
        12'h2de: data = 8'b00000000;	//         
        12'h2df: data = 8'b00000000;	//         

    // code xe2e (ฮ)
        12'h2e0: data = 8'b00000000;	//         
        12'h2e1: data = 8'b00000000;	//         
        12'h2e2: data = 8'b00000010;	//       * 
        12'h2e3: data = 8'b11111110;	// ******* 
        12'h2e4: data = 8'b00000010;	//       * 
        12'h2e5: data = 8'b00000010;	//       * 
        12'h2e6: data = 8'b11100010;	// ***   * 
        12'h2e7: data = 8'b11000010;	// **    * 
        12'h2e8: data = 8'b11000010;	// **    * 
        12'h2e9: data = 8'b00111100;	//   ****  
        12'h2ea: data = 8'b00000000;	//         
        12'h2eb: data = 8'b00000000;	//         
        12'h2ec: data = 8'b00000000;	//         
        12'h2ed: data = 8'b00000000;	//         
        12'h2ee: data = 8'b00000000;	//         
        12'h2ef: data = 8'b00000000;	//         

    // code xe2f (ฯ)
        12'h2f0: data = 8'b00000000;	//         
        12'h2f1: data = 8'b00000000;	//         
        12'h2f2: data = 8'b00000000;	//         
        12'h2f3: data = 8'b00100010;	//   *   * 
        12'h2f4: data = 8'b11000110;	// **   ** 
        12'h2f5: data = 8'b00110010;	//   **  * 
        12'h2f6: data = 8'b00110010;	//   **  * 
        12'h2f7: data = 8'b00000010;	//       * 
        12'h2f8: data = 8'b00000010;	//       * 
        12'h2f9: data = 8'b00011100;	//    ***  
        12'h2fa: data = 8'b00000000;	//         
        12'h2fb: data = 8'b00000000;	//         
        12'h2fc: data = 8'b00000000;	//         
        12'h2fd: data = 8'b00000000;	//         
        12'h2fe: data = 8'b00000000;	//         
        12'h2ff: data = 8'b00000000;	//         

    // code xe30 (ะ)
        12'h300: data = 8'b00000000;	//         
        12'h301: data = 8'b00000000;	//         
        12'h302: data = 8'b00000000;	//         
        12'h303: data = 8'b00000000;	//         
        12'h304: data = 8'b00000000;	//         
        12'h305: data = 8'b11000000;	// **      
        12'h306: data = 8'b11110000;	// ****    
        12'h307: data = 8'b00000000;	//         
        12'h308: data = 8'b11000000;	// **      
        12'h309: data = 8'b11110000;	// ****    
        12'h30a: data = 8'b00000000;	//         
        12'h30b: data = 8'b00000000;	//         
        12'h30c: data = 8'b00000000;	//         
        12'h30d: data = 8'b00000000;	//         
        12'h30e: data = 8'b00000000;	//         
        12'h30f: data = 8'b00000000;	//         

    // code xe31 (ั)
        12'h310: data = 8'b00000000;	//         
        12'h311: data = 8'b00000000;	//         
        12'h312: data = 8'b00000000;	//         
        12'h313: data = 8'b00000100;	//      *  
        12'h314: data = 8'b00000111;	//      ***
        12'h315: data = 8'b00000000;	//         
        12'h316: data = 8'b00000000;	//         
        12'h317: data = 8'b00000000;	//         
        12'h318: data = 8'b00000000;	//         
        12'h319: data = 8'b00000000;	//         
        12'h31a: data = 8'b00000000;	//         
        12'h31b: data = 8'b00000000;	//         
        12'h31c: data = 8'b00000000;	//         
        12'h31d: data = 8'b00000000;	//         
        12'h31e: data = 8'b00000000;	//         
        12'h31f: data = 8'b00000000;	//         

    // code xe32 (า)
        12'h320: data = 8'b00000000;	//         
        12'h321: data = 8'b00000000;	//         
        12'h322: data = 8'b00000000;	//         
        12'h323: data = 8'b11111000;	// *****   
        12'h324: data = 8'b00000100;	//      *  
        12'h325: data = 8'b00000100;	//      *  
        12'h326: data = 8'b00000100;	//      *  
        12'h327: data = 8'b00000100;	//      *  
        12'h328: data = 8'b00000100;	//      *  
        12'h329: data = 8'b00000100;	//      *  
        12'h32a: data = 8'b00000000;	//         
        12'h32b: data = 8'b00000000;	//         
        12'h32c: data = 8'b00000000;	//         
        12'h32d: data = 8'b00000000;	//         
        12'h32e: data = 8'b00000000;	//         
        12'h32f: data = 8'b00000000;	//         

    // code xe33 (ำ)
        12'h330: data = 8'b00000000;	//         
        12'h331: data = 8'b00000000;	//         
        12'h332: data = 8'b00000000;	//         
        12'h333: data = 8'b11111000;	// *****   
        12'h334: data = 8'b00000100;	//      *  
        12'h335: data = 8'b00000100;	//      *  
        12'h336: data = 8'b00000100;	//      *  
        12'h337: data = 8'b00000100;	//      *  
        12'h338: data = 8'b00000100;	//      *  
        12'h339: data = 8'b00000100;	//      *  
        12'h33a: data = 8'b00000000;	//         
        12'h33b: data = 8'b00000000;	//         
        12'h33c: data = 8'b00000000;	//         
        12'h33d: data = 8'b00000000;	//         
        12'h33e: data = 8'b00000000;	//         
        12'h33f: data = 8'b00000000;	//         

    // code xe34 (ิ)
        12'h340: data = 8'b00000000;	//         
        12'h341: data = 8'b00000000;	//         
        12'h342: data = 8'b00000000;	//         
        12'h343: data = 8'b00000000;	//         
        12'h344: data = 8'b00001111;	//     ****
        12'h345: data = 8'b00000000;	//         
        12'h346: data = 8'b00000000;	//         
        12'h347: data = 8'b00000000;	//         
        12'h348: data = 8'b00000000;	//         
        12'h349: data = 8'b00000000;	//         
        12'h34a: data = 8'b00000000;	//         
        12'h34b: data = 8'b00000000;	//         
        12'h34c: data = 8'b00000000;	//         
        12'h34d: data = 8'b00000000;	//         
        12'h34e: data = 8'b00000000;	//         
        12'h34f: data = 8'b00000000;	//         

    // code xe35 (ี)
        12'h350: data = 8'b00000000;	//         
        12'h351: data = 8'b00000000;	//         
        12'h352: data = 8'b00000000;	//         
        12'h353: data = 8'b00000001;	//        *
        12'h354: data = 8'b00001111;	//     ****
        12'h355: data = 8'b00000000;	//         
        12'h356: data = 8'b00000000;	//         
        12'h357: data = 8'b00000000;	//         
        12'h358: data = 8'b00000000;	//         
        12'h359: data = 8'b00000000;	//         
        12'h35a: data = 8'b00000000;	//         
        12'h35b: data = 8'b00000000;	//         
        12'h35c: data = 8'b00000000;	//         
        12'h35d: data = 8'b00000000;	//         
        12'h35e: data = 8'b00000000;	//         
        12'h35f: data = 8'b00000000;	//         

    // code xe36 (ึ)
        12'h360: data = 8'b00000000;	//         
        12'h361: data = 8'b00000000;	//         
        12'h362: data = 8'b00000000;	//         
        12'h363: data = 8'b00000011;	//       **
        12'h364: data = 8'b00001111;	//     ****
        12'h365: data = 8'b00000000;	//         
        12'h366: data = 8'b00000000;	//         
        12'h367: data = 8'b00000000;	//         
        12'h368: data = 8'b00000000;	//         
        12'h369: data = 8'b00000000;	//         
        12'h36a: data = 8'b00000000;	//         
        12'h36b: data = 8'b00000000;	//         
        12'h36c: data = 8'b00000000;	//         
        12'h36d: data = 8'b00000000;	//         
        12'h36e: data = 8'b00000000;	//         
        12'h36f: data = 8'b00000000;	//         

    // code xe37 (ื)
        12'h370: data = 8'b00000000;	//         
        12'h371: data = 8'b00000000;	//         
        12'h372: data = 8'b00000000;	//         
        12'h373: data = 8'b00000000;	//         
        12'h374: data = 8'b00001111;	//     ****
        12'h375: data = 8'b00000000;	//         
        12'h376: data = 8'b00000000;	//         
        12'h377: data = 8'b00000000;	//         
        12'h378: data = 8'b00000000;	//         
        12'h379: data = 8'b00000000;	//         
        12'h37a: data = 8'b00000000;	//         
        12'h37b: data = 8'b00000000;	//         
        12'h37c: data = 8'b00000000;	//         
        12'h37d: data = 8'b00000000;	//         
        12'h37e: data = 8'b00000000;	//         
        12'h37f: data = 8'b00000000;	//         

    // code xe38 (ุ)
        12'h380: data = 8'b00000000;	//         
        12'h381: data = 8'b00000000;	//         
        12'h382: data = 8'b00000000;	//         
        12'h383: data = 8'b00000000;	//         
        12'h384: data = 8'b00000000;	//         
        12'h385: data = 8'b00000000;	//         
        12'h386: data = 8'b00000000;	//         
        12'h387: data = 8'b00000000;	//         
        12'h388: data = 8'b00000000;	//         
        12'h389: data = 8'b00000000;	//         
        12'h38a: data = 8'b00000000;	//         
        12'h38b: data = 8'b00000001;	//        *
        12'h38c: data = 8'b00000001;	//        *
        12'h38d: data = 8'b00000000;	//         
        12'h38e: data = 8'b00000000;	//         
        12'h38f: data = 8'b00000000;	//         

    // code xe39 (ู)
        12'h390: data = 8'b00000000;	//         
        12'h391: data = 8'b00000000;	//         
        12'h392: data = 8'b00000000;	//         
        12'h393: data = 8'b00000000;	//         
        12'h394: data = 8'b00000000;	//         
        12'h395: data = 8'b00000000;	//         
        12'h396: data = 8'b00000000;	//         
        12'h397: data = 8'b00000000;	//         
        12'h398: data = 8'b00000000;	//         
        12'h399: data = 8'b00000000;	//         
        12'h39a: data = 8'b00000000;	//         
        12'h39b: data = 8'b00001001;	//     *  *
        12'h39c: data = 8'b00001111;	//     ****
        12'h39d: data = 8'b00000000;	//         
        12'h39e: data = 8'b00000000;	//         
        12'h39f: data = 8'b00000000;	//         

    // code xe40 (เ)
        12'h400: data = 8'b00000000;	//         
        12'h401: data = 8'b00000000;	//         
        12'h402: data = 8'b00000000;	//         
        12'h403: data = 8'b11000000;	// **      
        12'h404: data = 8'b11000000;	// **      
        12'h405: data = 8'b11000000;	// **      
        12'h406: data = 8'b11000000;	// **      
        12'h407: data = 8'b11000000;	// **      
        12'h408: data = 8'b11000000;	// **      
        12'h409: data = 8'b11000000;	// **      
        12'h40a: data = 8'b00000000;	//         
        12'h40b: data = 8'b00000000;	//         
        12'h40c: data = 8'b00000000;	//         
        12'h40d: data = 8'b00000000;	//         
        12'h40e: data = 8'b00000000;	//         
        12'h40f: data = 8'b00000000;	//         

    // code xe41 (แ)
        12'h410: data = 8'b00000000;	//         
        12'h411: data = 8'b00000000;	//         
        12'h412: data = 8'b00000000;	//         
        12'h413: data = 8'b11001000;	// **  *   
        12'h414: data = 8'b11001000;	// **  *   
        12'h415: data = 8'b11001000;	// **  *   
        12'h416: data = 8'b11001000;	// **  *   
        12'h417: data = 8'b11001000;	// **  *   
        12'h418: data = 8'b11001000;	// **  *   
        12'h419: data = 8'b11001000;	// **  *   
        12'h41a: data = 8'b00000000;	//         
        12'h41b: data = 8'b00000000;	//         
        12'h41c: data = 8'b00000000;	//         
        12'h41d: data = 8'b00000000;	//         
        12'h41e: data = 8'b00000000;	//         
        12'h41f: data = 8'b00000000;	//         

    // code xe42 (โ)
        12'h420: data = 8'b10000000;	// *       
        12'h421: data = 8'b11000000;	// **      
        12'h422: data = 8'b11000000;	// **      
        12'h423: data = 8'b11000000;	// **      
        12'h424: data = 8'b11000000;	// **      
        12'h425: data = 8'b11000000;	// **      
        12'h426: data = 8'b11000000;	// **      
        12'h427: data = 8'b11000000;	// **      
        12'h428: data = 8'b11000000;	// **      
        12'h429: data = 8'b11000000;	// **      
        12'h42a: data = 8'b00000000;	//         
        12'h42b: data = 8'b00000000;	//         
        12'h42c: data = 8'b00000000;	//         
        12'h42d: data = 8'b00000000;	//         
        12'h42e: data = 8'b00000000;	//         
        12'h42f: data = 8'b00000000;	//         

    // code xe43 (ใ)
        12'h430: data = 8'b11000000;	// **      
        12'h431: data = 8'b11000000;	// **      
        12'h432: data = 8'b11000000;	// **      
        12'h433: data = 8'b11000000;	// **      
        12'h434: data = 8'b11000000;	// **      
        12'h435: data = 8'b11000000;	// **      
        12'h436: data = 8'b11000000;	// **      
        12'h437: data = 8'b11000000;	// **      
        12'h438: data = 8'b11000000;	// **      
        12'h439: data = 8'b11000000;	// **      
        12'h43a: data = 8'b00000000;	//         
        12'h43b: data = 8'b00000000;	//         
        12'h43c: data = 8'b00000000;	//         
        12'h43d: data = 8'b00000000;	//         
        12'h43e: data = 8'b00000000;	//         
        12'h43f: data = 8'b00000000;	//         

    // code xe44 (ไ)
        12'h440: data = 8'b11000000;	// **      
        12'h441: data = 8'b11000000;	// **      
        12'h442: data = 8'b11000000;	// **      
        12'h443: data = 8'b11000000;	// **      
        12'h444: data = 8'b11000000;	// **      
        12'h445: data = 8'b11000000;	// **      
        12'h446: data = 8'b11000000;	// **      
        12'h447: data = 8'b11000000;	// **      
        12'h448: data = 8'b11000000;	// **      
        12'h449: data = 8'b11000000;	// **      
        12'h44a: data = 8'b00000000;	//         
        12'h44b: data = 8'b00000000;	//         
        12'h44c: data = 8'b00000000;	//         
        12'h44d: data = 8'b00000000;	//         
        12'h44e: data = 8'b00000000;	//         
        12'h44f: data = 8'b00000000;	//   

            default: data = 8'b00000000; // Default to zero
        endcase
 endmodule