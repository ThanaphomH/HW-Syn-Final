// *************************************************************
// Created by David J. Marion aka FPGA Dude
// A ROM containing patterns for ASCII values.
//
// Non-printable characters 00 - 1f, and 7f
// Printable characters 20 - 7e
//
// Not all character ROMs have been patterned.
// Only numbers, capital letters, some spec chars. 
//		Numbers       30 - 39
//   	Letters       41 - 5a 
//      (smiley face)   01
//		(space)         20
//		   .            2e
// 		   :            3a
//		   |	        7c	
//
// The 7-bit ASCII code for each character is used as
// the MSB of the address. The 4-bit LSB is the row value.
// *************************************************************

module ascii_rom(
        input clk, 
        input wire [10:0] addr,
        output reg [7:0] data
    );

    (* rom_style = "block" *) 

    reg [10:0] addr_reg;
    
    always @(posedge clk)
        addr_reg <= addr;
        
    always @*
        case(addr_reg)
    
    // code x41 (A)
        12'h410: data = 8'b00000000;	//         
        12'h411: data = 8'b00000000;	//         
        12'h412: data = 8'b00011000;	//    **   
        12'h413: data = 8'b00100100;	//   *  *  
        12'h414: data = 8'b11000010;	// **    * 
        12'h415: data = 8'b11000010;	// **    * 
        12'h416: data = 8'b11000010;	// **    * 
        12'h417: data = 8'b11111110;	// ******* 
        12'h418: data = 8'b11000010;	// **    * 
        12'h419: data = 8'b11000010;	// **    * 
        12'h41a: data = 8'b00000000;	//         
        12'h41b: data = 8'b00000000;	//         
        12'h41c: data = 8'b00000000;	//         
        12'h41d: data = 8'b00000000;	//         
        12'h41e: data = 8'b00000000;	//         
        12'h41f: data = 8'b00000000;	//         

    // code x42 (B)
        12'h420: data = 8'b00000000;	//         
        12'h421: data = 8'b00000000;	//         
        12'h422: data = 8'b11111100;	// ******  
        12'h423: data = 8'b11000010;	// **    * 
        12'h424: data = 8'b11000010;	// **    * 
        12'h425: data = 8'b11000000;	// **      
        12'h426: data = 8'b11111100;	// ******  
        12'h427: data = 8'b11000010;	// **    * 
        12'h428: data = 8'b11000010;	// **    * 
        12'h429: data = 8'b11111100;	// ******  
        12'h42a: data = 8'b00000000;	//         
        12'h42b: data = 8'b00000000;	//         
        12'h42c: data = 8'b00000000;	//         
        12'h42d: data = 8'b00000000;	//         
        12'h42e: data = 8'b00000000;	//         
        12'h42f: data = 8'b00000000;	//         

    // code x43 (C)
        12'h430: data = 8'b00000000;	//         
        12'h431: data = 8'b00000000;	//         
        12'h432: data = 8'b00111100;	//   ****  
        12'h433: data = 8'b00000010;	//       * 
        12'h434: data = 8'b11000010;	// **    * 
        12'h435: data = 8'b11000000;	// **      
        12'h436: data = 8'b11000000;	// **      
        12'h437: data = 8'b11000010;	// **    * 
        12'h438: data = 8'b11000010;	// **    * 
        12'h439: data = 8'b00111100;	//   ****  
        12'h43a: data = 8'b00000000;	//         
        12'h43b: data = 8'b00000000;	//         
        12'h43c: data = 8'b00000000;	//         
        12'h43d: data = 8'b00000000;	//         
        12'h43e: data = 8'b00000000;	//         
        12'h43f: data = 8'b00000000;	//         

    // code x44 (D)
        12'h440: data = 8'b00000000;	//         
        12'h441: data = 8'b00000000;	//         
        12'h442: data = 8'b11111000;	// *****   
        12'h443: data = 8'b11000100;	// **   *  
        12'h444: data = 8'b11000010;	// **    * 
        12'h445: data = 8'b11000010;	// **    * 
        12'h446: data = 8'b11000010;	// **    * 
        12'h447: data = 8'b11000010;	// **    * 
        12'h448: data = 8'b11000100;	// **   *  
        12'h449: data = 8'b11111000;	// *****   
        12'h44a: data = 8'b00000000;	//         
        12'h44b: data = 8'b00000000;	//         
        12'h44c: data = 8'b00000000;	//         
        12'h44d: data = 8'b00000000;	//         
        12'h44e: data = 8'b00000000;	//         
        12'h44f: data = 8'b00000000;	//         

    // code x45 (E)
        12'h450: data = 8'b00000000;	//         
        12'h451: data = 8'b00000000;	//         
        12'h452: data = 8'b11111100;	// ******  
        12'h453: data = 8'b11000000;	// **      
        12'h454: data = 8'b11000000;	// **      
        12'h455: data = 8'b11000000;	// **      
        12'h456: data = 8'b11111000;	// *****   
        12'h457: data = 8'b11000000;	// **      
        12'h458: data = 8'b11000000;	// **      
        12'h459: data = 8'b11111100;	// ******  
        12'h45a: data = 8'b00000000;	//         
        12'h45b: data = 8'b00000000;	//         
        12'h45c: data = 8'b00000000;	//         
        12'h45d: data = 8'b00000000;	//         
        12'h45e: data = 8'b00000000;	//         
        12'h45f: data = 8'b00000000;	//         

    // code x46 (F)
        12'h460: data = 8'b00000000;	//         
        12'h461: data = 8'b00000000;	//         
        12'h462: data = 8'b11111100;	// ******  
        12'h463: data = 8'b11000000;	// **      
        12'h464: data = 8'b11000000;	// **      
        12'h465: data = 8'b11000000;	// **      
        12'h466: data = 8'b11111000;	// *****   
        12'h467: data = 8'b11000000;	// **      
        12'h468: data = 8'b11000000;	// **      
        12'h469: data = 8'b11000000;	// **      
        12'h46a: data = 8'b00000000;	//         
        12'h46b: data = 8'b00000000;	//         
        12'h46c: data = 8'b00000000;	//         
        12'h46d: data = 8'b00000000;	//         
        12'h46e: data = 8'b00000000;	//         
        12'h46f: data = 8'b00000000;	//         

    // code x47 (G)
        12'h470: data = 8'b00000000;	//         
        12'h471: data = 8'b00000000;	//         
        12'h472: data = 8'b00111100;	//   ****  
        12'h473: data = 8'b00000010;	//       * 
        12'h474: data = 8'b11000000;	// **      
        12'h475: data = 8'b11000000;	// **      
        12'h476: data = 8'b11000110;	// **   ** 
        12'h477: data = 8'b11000010;	// **    * 
        12'h478: data = 8'b11000010;	// **    * 
        12'h479: data = 8'b00111100;	//   ****  
        12'h47a: data = 8'b00000000;	//         
        12'h47b: data = 8'b00000000;	//         
        12'h47c: data = 8'b00000000;	//         
        12'h47d: data = 8'b00000000;	//         
        12'h47e: data = 8'b00000000;	//         
        12'h47f: data = 8'b00000000;	//         

    // code x48 (H)
        12'h480: data = 8'b00000000;	//         
        12'h481: data = 8'b00000000;	//         
        12'h482: data = 8'b11000010;	// **    * 
        12'h483: data = 8'b11000010;	// **    * 
        12'h484: data = 8'b11000010;	// **    * 
        12'h485: data = 8'b11000010;	// **    * 
        12'h486: data = 8'b11111110;	// ******* 
        12'h487: data = 8'b11000010;	// **    * 
        12'h488: data = 8'b11000010;	// **    * 
        12'h489: data = 8'b11000010;	// **    * 
        12'h48a: data = 8'b00000000;	//         
        12'h48b: data = 8'b00000000;	//         
        12'h48c: data = 8'b00000000;	//         
        12'h48d: data = 8'b00000000;	//         
        12'h48e: data = 8'b00000000;	//         
        12'h48f: data = 8'b00000000;	//         

    // code x49 (I)
        12'h490: data = 8'b00000000;	//         
        12'h491: data = 8'b00000000;	//         
        12'h492: data = 8'b11000000;	// **      
        12'h493: data = 8'b11000000;	// **      
        12'h494: data = 8'b11000000;	// **      
        12'h495: data = 8'b11000000;	// **      
        12'h496: data = 8'b11000000;	// **      
        12'h497: data = 8'b11000000;	// **      
        12'h498: data = 8'b11000000;	// **      
        12'h499: data = 8'b11000000;	// **      
        12'h49a: data = 8'b00000000;	//         
        12'h49b: data = 8'b00000000;	//         
        12'h49c: data = 8'b00000000;	//         
        12'h49d: data = 8'b00000000;	//         
        12'h49e: data = 8'b00000000;	//         
        12'h49f: data = 8'b00000000;	//         

    // code x4a (J)
        12'h4a0: data = 8'b00000000;	//         
        12'h4a1: data = 8'b00000000;	//         
        12'h4a2: data = 8'b00010000;	//    *    
        12'h4a3: data = 8'b00010000;	//    *    
        12'h4a4: data = 8'b00010000;	//    *    
        12'h4a5: data = 8'b00010000;	//    *    
        12'h4a6: data = 8'b00010000;	//    *    
        12'h4a7: data = 8'b00010000;	//    *    
        12'h4a8: data = 8'b00010000;	//    *    
        12'h4a9: data = 8'b11100000;	// ***     
        12'h4aa: data = 8'b00000000;	//         
        12'h4ab: data = 8'b00000000;	//         
        12'h4ac: data = 8'b00000000;	//         
        12'h4ad: data = 8'b00000000;	//         
        12'h4ae: data = 8'b00000000;	//         
        12'h4af: data = 8'b00000000;	//         

    // code x4b (K)
        12'h4b0: data = 8'b00000000;	//         
        12'h4b1: data = 8'b00000000;	//         
        12'h4b2: data = 8'b11000010;	// **    * 
        12'h4b3: data = 8'b11000100;	// **   *  
        12'h4b4: data = 8'b11111000;	// *****   
        12'h4b5: data = 8'b11000100;	// **   *  
        12'h4b6: data = 8'b11000100;	// **   *  
        12'h4b7: data = 8'b11000010;	// **    * 
        12'h4b8: data = 8'b11000010;	// **    * 
        12'h4b9: data = 8'b11000010;	// **    * 
        12'h4ba: data = 8'b00000000;	//         
        12'h4bb: data = 8'b00000000;	//         
        12'h4bc: data = 8'b00000000;	//         
        12'h4bd: data = 8'b00000000;	//         
        12'h4be: data = 8'b00000000;	//         
        12'h4bf: data = 8'b00000000;	//         

    // code x4c (L)
        12'h4c0: data = 8'b00000000;	//         
        12'h4c1: data = 8'b00000000;	//         
        12'h4c2: data = 8'b11000000;	// **      
        12'h4c3: data = 8'b11000000;	// **      
        12'h4c4: data = 8'b11000000;	// **      
        12'h4c5: data = 8'b11000000;	// **      
        12'h4c6: data = 8'b11000000;	// **      
        12'h4c7: data = 8'b11000000;	// **      
        12'h4c8: data = 8'b11000000;	// **      
        12'h4c9: data = 8'b11111100;	// ******  
        12'h4ca: data = 8'b00000000;	//         
        12'h4cb: data = 8'b00000000;	//         
        12'h4cc: data = 8'b00000000;	//         
        12'h4cd: data = 8'b00000000;	//         
        12'h4ce: data = 8'b00000000;	//         
        12'h4cf: data = 8'b00000000;	//         

    // code x4d (M)
        12'h4d0: data = 8'b00000000;	//         
        12'h4d1: data = 8'b00000000;	//         
        12'h4d2: data = 8'b11100011;	// ***   **
        12'h4d3: data = 8'b11001001;	// **  *  *
        12'h4d4: data = 8'b11001001;	// **  *  *
        12'h4d5: data = 8'b11001001;	// **  *  *
        12'h4d6: data = 8'b11000001;	// **     *
        12'h4d7: data = 8'b11000001;	// **     *
        12'h4d8: data = 8'b11000001;	// **     *
        12'h4d9: data = 8'b11000001;	// **     *
        12'h4da: data = 8'b00000000;	//         
        12'h4db: data = 8'b00000000;	//         
        12'h4dc: data = 8'b00000000;	//         
        12'h4dd: data = 8'b00000000;	//         
        12'h4de: data = 8'b00000000;	//         
        12'h4df: data = 8'b00000000;	//         

    // code x4e (N)
        12'h4e0: data = 8'b00000000;	//         
        12'h4e1: data = 8'b00000000;	//         
        12'h4e2: data = 8'b11100010;	// ***   * 
        12'h4e3: data = 8'b11000010;	// **    * 
        12'h4e4: data = 8'b11000110;	// **   ** 
        12'h4e5: data = 8'b11000010;	// **    * 
        12'h4e6: data = 8'b11000010;	// **    * 
        12'h4e7: data = 8'b11000010;	// **    * 
        12'h4e8: data = 8'b11000010;	// **    * 
        12'h4e9: data = 8'b11000010;	// **    * 
        12'h4ea: data = 8'b00000000;	//         
        12'h4eb: data = 8'b00000000;	//         
        12'h4ec: data = 8'b00000000;	//         
        12'h4ed: data = 8'b00000000;	//         
        12'h4ee: data = 8'b00000000;	//         
        12'h4ef: data = 8'b00000000;	//         

    // code x4f (O)
        12'h4f0: data = 8'b00000000;	//         
        12'h4f1: data = 8'b00000000;	//         
        12'h4f2: data = 8'b00111100;	//   ****  
        12'h4f3: data = 8'b11000010;	// **    * 
        12'h4f4: data = 8'b11000010;	// **    * 
        12'h4f5: data = 8'b11000010;	// **    * 
        12'h4f6: data = 8'b11000010;	// **    * 
        12'h4f7: data = 8'b11000010;	// **    * 
        12'h4f8: data = 8'b11000010;	// **    * 
        12'h4f9: data = 8'b00111100;	//   ****  
        12'h4fa: data = 8'b00000000;	//         
        12'h4fb: data = 8'b00000000;	//         
        12'h4fc: data = 8'b00000000;	//         
        12'h4fd: data = 8'b00000000;	//         
        12'h4fe: data = 8'b00000000;	//         
        12'h4ff: data = 8'b00000000;	//         

    // code x50 (P)
        12'h500: data = 8'b00000000;	//         
        12'h501: data = 8'b00000000;	//         
        12'h502: data = 8'b11111100;	// ******  
        12'h503: data = 8'b11000010;	// **    * 
        12'h504: data = 8'b11000010;	// **    * 
        12'h505: data = 8'b11111100;	// ******  
        12'h506: data = 8'b11000000;	// **      
        12'h507: data = 8'b11000000;	// **      
        12'h508: data = 8'b11000000;	// **      
        12'h509: data = 8'b11000000;	// **      
        12'h50a: data = 8'b00000000;	//         
        12'h50b: data = 8'b00000000;	//         
        12'h50c: data = 8'b00000000;	//         
        12'h50d: data = 8'b00000000;	//         
        12'h50e: data = 8'b00000000;	//         
        12'h50f: data = 8'b00000000;	//         

    // code x51 (Q)
        12'h510: data = 8'b00000000;	//         
        12'h511: data = 8'b00000000;	//         
        12'h512: data = 8'b00111100;	//   ****  
        12'h513: data = 8'b11000010;	// **    * 
        12'h514: data = 8'b11000010;	// **    * 
        12'h515: data = 8'b11000010;	// **    * 
        12'h516: data = 8'b11000010;	// **    * 
        12'h517: data = 8'b11000010;	// **    * 
        12'h518: data = 8'b11000010;	// **    * 
        12'h519: data = 8'b00111100;	//   ****  
        12'h51a: data = 8'b00000000;	//         
        12'h51b: data = 8'b00000000;	//         
        12'h51c: data = 8'b00000000;	//         
        12'h51d: data = 8'b00000000;	//         
        12'h51e: data = 8'b00000000;	//         
        12'h51f: data = 8'b00000000;	//         

    // code x52 (R)
        12'h520: data = 8'b00000000;	//         
        12'h521: data = 8'b00000000;	//         
        12'h522: data = 8'b11111100;	// ******  
        12'h523: data = 8'b11000010;	// **    * 
        12'h524: data = 8'b11000010;	// **    * 
        12'h525: data = 8'b11000000;	// **      
        12'h526: data = 8'b11111100;	// ******  
        12'h527: data = 8'b11000010;	// **    * 
        12'h528: data = 8'b11000010;	// **    * 
        12'h529: data = 8'b11000010;	// **    * 
        12'h52a: data = 8'b00000000;	//         
        12'h52b: data = 8'b00000000;	//         
        12'h52c: data = 8'b00000000;	//         
        12'h52d: data = 8'b00000000;	//         
        12'h52e: data = 8'b00000000;	//         
        12'h52f: data = 8'b00000000;	//         

    // code x53 (S)
        12'h530: data = 8'b00000000;	//         
        12'h531: data = 8'b00000000;	//         
        12'h532: data = 8'b00111100;	//   ****  
        12'h533: data = 8'b11000010;	// **    * 
        12'h534: data = 8'b11000000;	// **      
        12'h535: data = 8'b00000000;	//         
        12'h536: data = 8'b00111100;	//   ****  
        12'h537: data = 8'b00000010;	//       * 
        12'h538: data = 8'b11000010;	// **    * 
        12'h539: data = 8'b00111100;	//   ****  
        12'h53a: data = 8'b00000000;	//         
        12'h53b: data = 8'b00000000;	//         
        12'h53c: data = 8'b00000000;	//         
        12'h53d: data = 8'b00000000;	//         
        12'h53e: data = 8'b00000000;	//         
        12'h53f: data = 8'b00000000;	//         

    // code x54 (T)
        12'h540: data = 8'b00000000;	//         
        12'h541: data = 8'b00000000;	//         
        12'h542: data = 8'b11111100;	// ******  
        12'h543: data = 8'b00010000;	//    *    
        12'h544: data = 8'b00010000;	//    *    
        12'h545: data = 8'b00010000;	//    *    
        12'h546: data = 8'b00010000;	//    *    
        12'h547: data = 8'b00010000;	//    *    
        12'h548: data = 8'b00010000;	//    *    
        12'h549: data = 8'b00010000;	//    *    
        12'h54a: data = 8'b00000000;	//         
        12'h54b: data = 8'b00000000;	//         
        12'h54c: data = 8'b00000000;	//         
        12'h54d: data = 8'b00000000;	//         
        12'h54e: data = 8'b00000000;	//         
        12'h54f: data = 8'b00000000;	//         

    // code x55 (U)
        12'h550: data = 8'b00000000;	//         
        12'h551: data = 8'b00000000;	//         
        12'h552: data = 8'b11000010;	// **    * 
        12'h553: data = 8'b11000010;	// **    * 
        12'h554: data = 8'b11000010;	// **    * 
        12'h555: data = 8'b11000010;	// **    * 
        12'h556: data = 8'b11000010;	// **    * 
        12'h557: data = 8'b11000010;	// **    * 
        12'h558: data = 8'b11000010;	// **    * 
        12'h559: data = 8'b00111100;	//   ****  
        12'h55a: data = 8'b00000000;	//         
        12'h55b: data = 8'b00000000;	//         
        12'h55c: data = 8'b00000000;	//         
        12'h55d: data = 8'b00000000;	//         
        12'h55e: data = 8'b00000000;	//         
        12'h55f: data = 8'b00000000;	//         

    // code x56 (V)
        12'h560: data = 8'b00000000;	//         
        12'h561: data = 8'b00000000;	//         
        12'h562: data = 8'b11000010;	// **    * 
        12'h563: data = 8'b11000010;	// **    * 
        12'h564: data = 8'b11000010;	// **    * 
        12'h565: data = 8'b11000010;	// **    * 
        12'h566: data = 8'b11000010;	// **    * 
        12'h567: data = 8'b11000010;	// **    * 
        12'h568: data = 8'b00100100;	//   *  *  
        12'h569: data = 8'b00011000;	//    **   
        12'h56a: data = 8'b00000000;	//         
        12'h56b: data = 8'b00000000;	//         
        12'h56c: data = 8'b00000000;	//         
        12'h56d: data = 8'b00000000;	//         
        12'h56e: data = 8'b00000000;	//         
        12'h56f: data = 8'b00000000;	//         

    // code x57 (W)
        12'h570: data = 8'b00000000;	//         
        12'h571: data = 8'b00000000;	//         
        12'h572: data = 8'b11000001;	// **     *
        12'h573: data = 8'b11000001;	// **     *
        12'h574: data = 8'b11000001;	// **     *
        12'h575: data = 8'b11001001;	// **  *  *
        12'h576: data = 8'b11001001;	// **  *  *
        12'h577: data = 8'b11001001;	// **  *  *
        12'h578: data = 8'b11001001;	// **  *  *
        12'h579: data = 8'b00100010;	//   *   * 
        12'h57a: data = 8'b00000000;	//         
        12'h57b: data = 8'b00000000;	//         
        12'h57c: data = 8'b00000000;	//         
        12'h57d: data = 8'b00000000;	//         
        12'h57e: data = 8'b00000000;	//         
        12'h57f: data = 8'b00000000;	//         

    // code x58 (X)
        12'h580: data = 8'b00000000;	//         
        12'h581: data = 8'b00000000;	//         
        12'h582: data = 8'b00000100;	//      *  
        12'h583: data = 8'b11000100;	// **   *  
        12'h584: data = 8'b00000000;	//         
        12'h585: data = 8'b00010000;	//    *    
        12'h586: data = 8'b00010000;	//    *    
        12'h587: data = 8'b00000000;	//         
        12'h588: data = 8'b11000100;	// **   *  
        12'h589: data = 8'b11000100;	// **   *  
        12'h58a: data = 8'b00000000;	//         
        12'h58b: data = 8'b00000000;	//         
        12'h58c: data = 8'b00000000;	//         
        12'h58d: data = 8'b00000000;	//         
        12'h58e: data = 8'b00000000;	//         
        12'h58f: data = 8'b00000000;	//         

    // code x59 (Y)
        12'h590: data = 8'b00000000;	//         
        12'h591: data = 8'b00000000;	//         
        12'h592: data = 8'b11000100;	// **   *  
        12'h593: data = 8'b11000100;	// **   *  
        12'h594: data = 8'b11000100;	// **   *  
        12'h595: data = 8'b00111000;	//   ***   
        12'h596: data = 8'b00010000;	//    *    
        12'h597: data = 8'b00010000;	//    *    
        12'h598: data = 8'b00010000;	//    *    
        12'h599: data = 8'b00010000;	//    *    
        12'h59a: data = 8'b00000000;	//         
        12'h59b: data = 8'b00000000;	//         
        12'h59c: data = 8'b00000000;	//         
        12'h59d: data = 8'b00000000;	//         
        12'h59e: data = 8'b00000000;	//         
        12'h59f: data = 8'b00000000;	//         

    // code x5a (Z)
        12'h5a0: data = 8'b00000000;	//         
        12'h5a1: data = 8'b00000000;	//         
        12'h5a2: data = 8'b11111100;	// ******  
        12'h5a3: data = 8'b00000100;	//      *  
        12'h5a4: data = 8'b00001000;	//     *   
        12'h5a5: data = 8'b00001000;	//     *   
        12'h5a6: data = 8'b00010000;	//    *    
        12'h5a7: data = 8'b00100000;	//   *     
        12'h5a8: data = 8'b11000000;	// **      
        12'h5a9: data = 8'b11111100;	// ******  
        12'h5aa: data = 8'b00000000;	//         
        12'h5ab: data = 8'b00000000;	//         
        12'h5ac: data = 8'b00000000;	//         
        12'h5ad: data = 8'b00000000;	//         
        12'h5ae: data = 8'b00000000;	//         
        12'h5af: data = 8'b00000000;	//         

    // code x61 (a)
        12'h610: data = 8'b00000000;	//         
        12'h611: data = 8'b00000000;	//         
        12'h612: data = 8'b00000000;	//         
        12'h613: data = 8'b00111100;	//   ****  
        12'h614: data = 8'b00000010;	//       * 
        12'h615: data = 8'b00000010;	//       * 
        12'h616: data = 8'b00111110;	//   ***** 
        12'h617: data = 8'b11000010;	// **    * 
        12'h618: data = 8'b11000010;	// **    * 
        12'h619: data = 8'b00111110;	//   ***** 
        12'h61a: data = 8'b00000000;	//         
        12'h61b: data = 8'b00000000;	//         
        12'h61c: data = 8'b00000000;	//         
        12'h61d: data = 8'b00000000;	//         
        12'h61e: data = 8'b00000000;	//         
        12'h61f: data = 8'b00000000;	//         

    // code x62 (b)
        12'h620: data = 8'b00000000;	//         
        12'h621: data = 8'b11000000;	// **      
        12'h622: data = 8'b11000000;	// **      
        12'h623: data = 8'b11111100;	// ******  
        12'h624: data = 8'b11000010;	// **    * 
        12'h625: data = 8'b11000010;	// **    * 
        12'h626: data = 8'b11000010;	// **    * 
        12'h627: data = 8'b11000010;	// **    * 
        12'h628: data = 8'b11000010;	// **    * 
        12'h629: data = 8'b11111100;	// ******  
        12'h62a: data = 8'b00000000;	//         
        12'h62b: data = 8'b00000000;	//         
        12'h62c: data = 8'b00000000;	//         
        12'h62d: data = 8'b00000000;	//         
        12'h62e: data = 8'b00000000;	//         
        12'h62f: data = 8'b00000000;	//         

    // code x63 (c)
        12'h630: data = 8'b00000000;	//         
        12'h631: data = 8'b00000000;	//         
        12'h632: data = 8'b00000000;	//         
        12'h633: data = 8'b00111100;	//   ****  
        12'h634: data = 8'b11000000;	// **      
        12'h635: data = 8'b11000010;	// **    * 
        12'h636: data = 8'b11000000;	// **      
        12'h637: data = 8'b11000000;	// **      
        12'h638: data = 8'b11000010;	// **    * 
        12'h639: data = 8'b00111100;	//   ****  
        12'h63a: data = 8'b00000000;	//         
        12'h63b: data = 8'b00000000;	//         
        12'h63c: data = 8'b00000000;	//         
        12'h63d: data = 8'b00000000;	//         
        12'h63e: data = 8'b00000000;	//         
        12'h63f: data = 8'b00000000;	//         

    // code x64 (d)
        12'h640: data = 8'b00000000;	//         
        12'h641: data = 8'b00000010;	//       * 
        12'h642: data = 8'b00000010;	//       * 
        12'h643: data = 8'b00111110;	//   ***** 
        12'h644: data = 8'b11000010;	// **    * 
        12'h645: data = 8'b11000010;	// **    * 
        12'h646: data = 8'b11000010;	// **    * 
        12'h647: data = 8'b11000010;	// **    * 
        12'h648: data = 8'b11000010;	// **    * 
        12'h649: data = 8'b00111110;	//   ***** 
        12'h64a: data = 8'b00000000;	//         
        12'h64b: data = 8'b00000000;	//         
        12'h64c: data = 8'b00000000;	//         
        12'h64d: data = 8'b00000000;	//         
        12'h64e: data = 8'b00000000;	//         
        12'h64f: data = 8'b00000000;	//         

    // code x65 (e)
        12'h650: data = 8'b00000000;	//         
        12'h651: data = 8'b00000000;	//         
        12'h652: data = 8'b00000000;	//         
        12'h653: data = 8'b00111100;	//   ****  
        12'h654: data = 8'b11000000;	// **      
        12'h655: data = 8'b11000010;	// **    * 
        12'h656: data = 8'b11000010;	// **    * 
        12'h657: data = 8'b11111100;	// ******  
        12'h658: data = 8'b11000000;	// **      
        12'h659: data = 8'b00111100;	//   ****  
        12'h65a: data = 8'b00000000;	//         
        12'h65b: data = 8'b00000000;	//         
        12'h65c: data = 8'b00000000;	//         
        12'h65d: data = 8'b00000000;	//         
        12'h65e: data = 8'b00000000;	//         
        12'h65f: data = 8'b00000000;	//         

    // code x66 (f)
        12'h660: data = 8'b00000000;	//         
        12'h661: data = 8'b00110000;	//   **    
        12'h662: data = 8'b11000000;	// **      
        12'h663: data = 8'b11000000;	// **      
        12'h664: data = 8'b11000000;	// **      
        12'h665: data = 8'b11110000;	// ****    
        12'h666: data = 8'b11000000;	// **      
        12'h667: data = 8'b11000000;	// **      
        12'h668: data = 8'b11000000;	// **      
        12'h669: data = 8'b11000000;	// **      
        12'h66a: data = 8'b00000000;	//         
        12'h66b: data = 8'b00000000;	//         
        12'h66c: data = 8'b00000000;	//         
        12'h66d: data = 8'b00000000;	//         
        12'h66e: data = 8'b00000000;	//         
        12'h66f: data = 8'b00000000;	//         

    // code x67 (g)
        12'h670: data = 8'b00000000;	//         
        12'h671: data = 8'b00000000;	//         
        12'h672: data = 8'b00000100;	//      *  
        12'h673: data = 8'b00111110;	//   ***** 
        12'h674: data = 8'b11000010;	// **    * 
        12'h675: data = 8'b11000010;	// **    * 
        12'h676: data = 8'b00000000;	//         
        12'h677: data = 8'b00111100;	//   ****  
        12'h678: data = 8'b00001000;	//     *   
        12'h679: data = 8'b00111100;	//   ****  
        12'h67a: data = 8'b11000010;	// **    * 
        12'h67b: data = 8'b11000010;	// **    * 
        12'h67c: data = 8'b00000000;	//         
        12'h67d: data = 8'b00000000;	//         
        12'h67e: data = 8'b00000000;	//         
        12'h67f: data = 8'b00000000;	//         

    // code x68 (h)
        12'h680: data = 8'b00000000;	//         
        12'h681: data = 8'b11000000;	// **      
        12'h682: data = 8'b11000000;	// **      
        12'h683: data = 8'b11111100;	// ******  
        12'h684: data = 8'b11000010;	// **    * 
        12'h685: data = 8'b11000010;	// **    * 
        12'h686: data = 8'b11000010;	// **    * 
        12'h687: data = 8'b11000010;	// **    * 
        12'h688: data = 8'b11000010;	// **    * 
        12'h689: data = 8'b11000010;	// **    * 
        12'h68a: data = 8'b00000000;	//         
        12'h68b: data = 8'b00000000;	//         
        12'h68c: data = 8'b00000000;	//         
        12'h68d: data = 8'b00000000;	//         
        12'h68e: data = 8'b00000000;	//         
        12'h68f: data = 8'b00000000;	//         

    // code x69 (i)
        12'h690: data = 8'b00000000;	//         
        12'h691: data = 8'b11000000;	// **      
        12'h692: data = 8'b00000000;	//         
        12'h693: data = 8'b00000000;	//         
        12'h694: data = 8'b11000000;	// **      
        12'h695: data = 8'b11000000;	// **      
        12'h696: data = 8'b11000000;	// **      
        12'h697: data = 8'b11000000;	// **      
        12'h698: data = 8'b11000000;	// **      
        12'h699: data = 8'b11000000;	// **      
        12'h69a: data = 8'b00000000;	//         
        12'h69b: data = 8'b00000000;	//         
        12'h69c: data = 8'b00000000;	//         
        12'h69d: data = 8'b00000000;	//         
        12'h69e: data = 8'b00000000;	//         
        12'h69f: data = 8'b00000000;	//         

    // code x6a (j)
        12'h6a0: data = 8'b00000000;	//         
        12'h6a1: data = 8'b11000000;	// **      
        12'h6a2: data = 8'b00000000;	//         
        12'h6a3: data = 8'b00000000;	//         
        12'h6a4: data = 8'b11000000;	// **      
        12'h6a5: data = 8'b11000000;	// **      
        12'h6a6: data = 8'b11000000;	// **      
        12'h6a7: data = 8'b11000000;	// **      
        12'h6a8: data = 8'b11000000;	// **      
        12'h6a9: data = 8'b11000000;	// **      
        12'h6aa: data = 8'b11000000;	// **      
        12'h6ab: data = 8'b10000000;	// *       
        12'h6ac: data = 8'b00000000;	//         
        12'h6ad: data = 8'b00000000;	//         
        12'h6ae: data = 8'b00000000;	//         
        12'h6af: data = 8'b00000000;	//         

    // code x6b (k)
        12'h6b0: data = 8'b00000000;	//         
        12'h6b1: data = 8'b11000000;	// **      
        12'h6b2: data = 8'b11000000;	// **      
        12'h6b3: data = 8'b11000100;	// **   *  
        12'h6b4: data = 8'b11001000;	// **  *   
        12'h6b5: data = 8'b11000000;	// **      
        12'h6b6: data = 8'b11110000;	// ****    
        12'h6b7: data = 8'b11001000;	// **  *   
        12'h6b8: data = 8'b11000100;	// **   *  
        12'h6b9: data = 8'b11000100;	// **   *  
        12'h6ba: data = 8'b00000000;	//         
        12'h6bb: data = 8'b00000000;	//         
        12'h6bc: data = 8'b00000000;	//         
        12'h6bd: data = 8'b00000000;	//         
        12'h6be: data = 8'b00000000;	//         
        12'h6bf: data = 8'b00000000;	//         

    // code x6c (l)
        12'h6c0: data = 8'b00000000;	//         
        12'h6c1: data = 8'b11000000;	// **      
        12'h6c2: data = 8'b11000000;	// **      
        12'h6c3: data = 8'b11000000;	// **      
        12'h6c4: data = 8'b11000000;	// **      
        12'h6c5: data = 8'b11000000;	// **      
        12'h6c6: data = 8'b11000000;	// **      
        12'h6c7: data = 8'b11000000;	// **      
        12'h6c8: data = 8'b11000000;	// **      
        12'h6c9: data = 8'b11000000;	// **      
        12'h6ca: data = 8'b00000000;	//         
        12'h6cb: data = 8'b00000000;	//         
        12'h6cc: data = 8'b00000000;	//         
        12'h6cd: data = 8'b00000000;	//         
        12'h6ce: data = 8'b00000000;	//         
        12'h6cf: data = 8'b00000000;	//         

    // code x6d (m)
        12'h6d0: data = 8'b00000000;	//         
        12'h6d1: data = 8'b00000000;	//         
        12'h6d2: data = 8'b00000000;	//         
        12'h6d3: data = 8'b11100010;	// ***   * 
        12'h6d4: data = 8'b11001001;	// **  *  *
        12'h6d5: data = 8'b11001001;	// **  *  *
        12'h6d6: data = 8'b11001001;	// **  *  *
        12'h6d7: data = 8'b11001001;	// **  *  *
        12'h6d8: data = 8'b11001001;	// **  *  *
        12'h6d9: data = 8'b11001001;	// **  *  *
        12'h6da: data = 8'b00000000;	//         
        12'h6db: data = 8'b00000000;	//         
        12'h6dc: data = 8'b00000000;	//         
        12'h6dd: data = 8'b00000000;	//         
        12'h6de: data = 8'b00000000;	//         
        12'h6df: data = 8'b00000000;	//         

    // code x6e (n)
        12'h6e0: data = 8'b00000000;	//         
        12'h6e1: data = 8'b00000000;	//         
        12'h6e2: data = 8'b00000000;	//         
        12'h6e3: data = 8'b11111100;	// ******  
        12'h6e4: data = 8'b11000010;	// **    * 
        12'h6e5: data = 8'b11000010;	// **    * 
        12'h6e6: data = 8'b11000010;	// **    * 
        12'h6e7: data = 8'b11000010;	// **    * 
        12'h6e8: data = 8'b11000010;	// **    * 
        12'h6e9: data = 8'b11000010;	// **    * 
        12'h6ea: data = 8'b00000000;	//         
        12'h6eb: data = 8'b00000000;	//         
        12'h6ec: data = 8'b00000000;	//         
        12'h6ed: data = 8'b00000000;	//         
        12'h6ee: data = 8'b00000000;	//         
        12'h6ef: data = 8'b00000000;	//         

    // code x6f (o)
        12'h6f0: data = 8'b00000000;	//         
        12'h6f1: data = 8'b00000000;	//         
        12'h6f2: data = 8'b00000000;	//         
        12'h6f3: data = 8'b00111100;	//   ****  
        12'h6f4: data = 8'b11000010;	// **    * 
        12'h6f5: data = 8'b11000010;	// **    * 
        12'h6f6: data = 8'b11000010;	// **    * 
        12'h6f7: data = 8'b11000010;	// **    * 
        12'h6f8: data = 8'b11000010;	// **    * 
        12'h6f9: data = 8'b00111100;	//   ****  
        12'h6fa: data = 8'b00000000;	//         
        12'h6fb: data = 8'b00000000;	//         
        12'h6fc: data = 8'b00000000;	//         
        12'h6fd: data = 8'b00000000;	//         
        12'h6fe: data = 8'b00000000;	//         
        12'h6ff: data = 8'b00000000;	//         

    // code x70 (p)
        12'h700: data = 8'b00000000;	//         
        12'h701: data = 8'b00000000;	//         
        12'h702: data = 8'b00000000;	//         
        12'h703: data = 8'b11111100;	// ******  
        12'h704: data = 8'b11000010;	// **    * 
        12'h705: data = 8'b11000010;	// **    * 
        12'h706: data = 8'b11000010;	// **    * 
        12'h707: data = 8'b11000010;	// **    * 
        12'h708: data = 8'b11000010;	// **    * 
        12'h709: data = 8'b11111100;	// ******  
        12'h70a: data = 8'b11000000;	// **      
        12'h70b: data = 8'b11000000;	// **      
        12'h70c: data = 8'b00000000;	//         
        12'h70d: data = 8'b00000000;	//         
        12'h70e: data = 8'b00000000;	//         
        12'h70f: data = 8'b00000000;	//         

    // code x71 (q)
        12'h710: data = 8'b00000000;	//         
        12'h711: data = 8'b00000000;	//         
        12'h712: data = 8'b00000000;	//         
        12'h713: data = 8'b00111110;	//   ***** 
        12'h714: data = 8'b11000010;	// **    * 
        12'h715: data = 8'b11000010;	// **    * 
        12'h716: data = 8'b11000010;	// **    * 
        12'h717: data = 8'b11000010;	// **    * 
        12'h718: data = 8'b11000010;	// **    * 
        12'h719: data = 8'b00111110;	//   ***** 
        12'h71a: data = 8'b00000010;	//       * 
        12'h71b: data = 8'b00000010;	//       * 
        12'h71c: data = 8'b00000000;	//         
        12'h71d: data = 8'b00000000;	//         
        12'h71e: data = 8'b00000000;	//         
        12'h71f: data = 8'b00000000;	//         

    // code x72 (r)
        12'h720: data = 8'b00000000;	//         
        12'h721: data = 8'b00000000;	//         
        12'h722: data = 8'b00000000;	//         
        12'h723: data = 8'b11111000;	// *****   
        12'h724: data = 8'b11000100;	// **   *  
        12'h725: data = 8'b11000000;	// **      
        12'h726: data = 8'b11000000;	// **      
        12'h727: data = 8'b11000000;	// **      
        12'h728: data = 8'b11000000;	// **      
        12'h729: data = 8'b11000000;	// **      
        12'h72a: data = 8'b00000000;	//         
        12'h72b: data = 8'b00000000;	//         
        12'h72c: data = 8'b00000000;	//         
        12'h72d: data = 8'b00000000;	//         
        12'h72e: data = 8'b00000000;	//         
        12'h72f: data = 8'b00000000;	//         

    // code x73 (s)
        12'h730: data = 8'b00000000;	//         
        12'h731: data = 8'b00000000;	//         
        12'h732: data = 8'b00000000;	//         
        12'h733: data = 8'b00111100;	//   ****  
        12'h734: data = 8'b11000000;	// **      
        12'h735: data = 8'b00000000;	//         
        12'h736: data = 8'b00111000;	//   ***   
        12'h737: data = 8'b00000100;	//      *  
        12'h738: data = 8'b00000100;	//      *  
        12'h739: data = 8'b11111000;	// *****   
        12'h73a: data = 8'b00000000;	//         
        12'h73b: data = 8'b00000000;	//         
        12'h73c: data = 8'b00000000;	//         
        12'h73d: data = 8'b00000000;	//         
        12'h73e: data = 8'b00000000;	//         
        12'h73f: data = 8'b00000000;	//         

    // code x74 (t)
        12'h740: data = 8'b00000000;	//         
        12'h741: data = 8'b00100000;	//   *     
        12'h742: data = 8'b00100000;	//   *     
        12'h743: data = 8'b11110000;	// ****    
        12'h744: data = 8'b00100000;	//   *     
        12'h745: data = 8'b00100000;	//   *     
        12'h746: data = 8'b00100000;	//   *     
        12'h747: data = 8'b00100000;	//   *     
        12'h748: data = 8'b00100000;	//   *     
        12'h749: data = 8'b00010000;	//    *    
        12'h74a: data = 8'b00000000;	//         
        12'h74b: data = 8'b00000000;	//         
        12'h74c: data = 8'b00000000;	//         
        12'h74d: data = 8'b00000000;	//         
        12'h74e: data = 8'b00000000;	//         
        12'h74f: data = 8'b00000000;	//         

    // code x75 (u)
        12'h750: data = 8'b00000000;	//         
        12'h751: data = 8'b00000000;	//         
        12'h752: data = 8'b00000000;	//         
        12'h753: data = 8'b11000010;	// **    * 
        12'h754: data = 8'b11000010;	// **    * 
        12'h755: data = 8'b11000010;	// **    * 
        12'h756: data = 8'b11000010;	// **    * 
        12'h757: data = 8'b11000010;	// **    * 
        12'h758: data = 8'b11000010;	// **    * 
        12'h759: data = 8'b00111110;	//   ***** 
        12'h75a: data = 8'b00000000;	//         
        12'h75b: data = 8'b00000000;	//         
        12'h75c: data = 8'b00000000;	//         
        12'h75d: data = 8'b00000000;	//         
        12'h75e: data = 8'b00000000;	//         
        12'h75f: data = 8'b00000000;	//         

    // code x76 (v)
        12'h760: data = 8'b00000000;	//         
        12'h761: data = 8'b00000000;	//         
        12'h762: data = 8'b00000000;	//         
        12'h763: data = 8'b11000010;	// **    * 
        12'h764: data = 8'b11000010;	// **    * 
        12'h765: data = 8'b11000010;	// **    * 
        12'h766: data = 8'b11000010;	// **    * 
        12'h767: data = 8'b11000010;	// **    * 
        12'h768: data = 8'b00100100;	//   *  *  
        12'h769: data = 8'b00011000;	//    **   
        12'h76a: data = 8'b00000000;	//         
        12'h76b: data = 8'b00000000;	//         
        12'h76c: data = 8'b00000000;	//         
        12'h76d: data = 8'b00000000;	//         
        12'h76e: data = 8'b00000000;	//         
        12'h76f: data = 8'b00000000;	//         

    // code x77 (w)
        12'h770: data = 8'b00000000;	//         
        12'h771: data = 8'b00000000;	//         
        12'h772: data = 8'b00000000;	//         
        12'h773: data = 8'b11000010;	// **    * 
        12'h774: data = 8'b11000010;	// **    * 
        12'h775: data = 8'b11000010;	// **    * 
        12'h776: data = 8'b11000010;	// **    * 
        12'h777: data = 8'b11000010;	// **    * 
        12'h778: data = 8'b11000010;	// **    * 
        12'h779: data = 8'b00100100;	//   *  *  
        12'h77a: data = 8'b00000000;	//         
        12'h77b: data = 8'b00000000;	//         
        12'h77c: data = 8'b00000000;	//         
        12'h77d: data = 8'b00000000;	//         
        12'h77e: data = 8'b00000000;	//         
        12'h77f: data = 8'b00000000;	//         

    // code x78 (x)
        12'h780: data = 8'b00000000;	//         
        12'h781: data = 8'b00000000;	//         
        12'h782: data = 8'b00000000;	//         
        12'h783: data = 8'b11000000;	// **      
        12'h784: data = 8'b00100100;	//   *  *  
        12'h785: data = 8'b00000000;	//         
        12'h786: data = 8'b00011000;	//    **   
        12'h787: data = 8'b00100100;	//   *  *  
        12'h788: data = 8'b11000010;	// **    * 
        12'h789: data = 8'b11000010;	// **    * 
        12'h78a: data = 8'b00000000;	//         
        12'h78b: data = 8'b00000000;	//         
        12'h78c: data = 8'b00000000;	//         
        12'h78d: data = 8'b00000000;	//         
        12'h78e: data = 8'b00000000;	//         
        12'h78f: data = 8'b00000000;	//         

    // code x79 (y)
        12'h790: data = 8'b00000000;	//         
        12'h791: data = 8'b00000000;	//         
        12'h792: data = 8'b00000000;	//         
        12'h793: data = 8'b11000010;	// **    * 
        12'h794: data = 8'b11000010;	// **    * 
        12'h795: data = 8'b11000010;	// **    * 
        12'h796: data = 8'b11000010;	// **    * 
        12'h797: data = 8'b11000010;	// **    * 
        12'h798: data = 8'b11000010;	// **    * 
        12'h799: data = 8'b00111110;	//   ***** 
        12'h79a: data = 8'b00000010;	//       * 
        12'h79b: data = 8'b00111100;	//   ****  
        12'h79c: data = 8'b00000000;	//         
        12'h79d: data = 8'b00000000;	//         
        12'h79e: data = 8'b00000000;	//         
        12'h79f: data = 8'b00000000;	//         

    // code x7a (z)
        12'h7a0: data = 8'b00000000;	//         
        12'h7a1: data = 8'b00000000;	//         
        12'h7a2: data = 8'b00000000;	//         
        12'h7a3: data = 8'b00000000;	//         
        12'h7a4: data = 8'b00001000;	//     *   
        12'h7a5: data = 8'b00010000;	//    *    
        12'h7a6: data = 8'b00010000;	//    *    
        12'h7a7: data = 8'b01000000;	//  *      
        12'h7a8: data = 8'b11000000;	// **      
        12'h7a9: data = 8'b11111000;	// *****   
        12'h7aa: data = 8'b00000000;	//         
        12'h7ab: data = 8'b00000000;	//         
        12'h7ac: data = 8'b00000000;	//         
        12'h7ad: data = 8'b00000000;	//         
        12'h7ae: data = 8'b00000000;	//         
        12'h7af: data = 8'b00000000;	//         

    // code x30 (0)
        12'h300: data = 8'b00000000;	//         
        12'h301: data = 8'b00000000;	//         
        12'h302: data = 8'b00111100;	//   ****  
        12'h303: data = 8'b11000010;	// **    * 
        12'h304: data = 8'b11000010;	// **    * 
        12'h305: data = 8'b11000010;	// **    * 
        12'h306: data = 8'b11000110;	// **   ** 
        12'h307: data = 8'b11000010;	// **    * 
        12'h308: data = 8'b11100010;	// ***   * 
        12'h309: data = 8'b00111100;	//   ****  
        12'h30a: data = 8'b00000000;	//         
        12'h30b: data = 8'b00000000;	//         
        12'h30c: data = 8'b00000000;	//         
        12'h30d: data = 8'b00000000;	//         
        12'h30e: data = 8'b00000000;	//         
        12'h30f: data = 8'b00000000;	//         

    // code x31 (1)
        12'h310: data = 8'b00000000;	//         
        12'h311: data = 8'b00000000;	//         
        12'h312: data = 8'b00100000;	//   *     
        12'h313: data = 8'b11100000;	// ***     
        12'h314: data = 8'b00100000;	//   *     
        12'h315: data = 8'b00100000;	//   *     
        12'h316: data = 8'b00100000;	//   *     
        12'h317: data = 8'b00100000;	//   *     
        12'h318: data = 8'b00100000;	//   *     
        12'h319: data = 8'b11110000;	// ****    
        12'h31a: data = 8'b00000000;	//         
        12'h31b: data = 8'b00000000;	//         
        12'h31c: data = 8'b00000000;	//         
        12'h31d: data = 8'b00000000;	//         
        12'h31e: data = 8'b00000000;	//         
        12'h31f: data = 8'b00000000;	//         

    // code x32 (2)
        12'h320: data = 8'b00000000;	//         
        12'h321: data = 8'b00000000;	//         
        12'h322: data = 8'b00111100;	//   ****  
        12'h323: data = 8'b11000010;	// **    * 
        12'h324: data = 8'b00000010;	//       * 
        12'h325: data = 8'b00000010;	//       * 
        12'h326: data = 8'b00011100;	//    ***  
        12'h327: data = 8'b00100000;	//   *     
        12'h328: data = 8'b11000000;	// **      
        12'h329: data = 8'b11111110;	// ******* 
        12'h32a: data = 8'b00000000;	//         
        12'h32b: data = 8'b00000000;	//         
        12'h32c: data = 8'b00000000;	//         
        12'h32d: data = 8'b00000000;	//         
        12'h32e: data = 8'b00000000;	//         
        12'h32f: data = 8'b00000000;	//         

    // code x33 (3)
        12'h330: data = 8'b00000000;	//         
        12'h331: data = 8'b00000000;	//         
        12'h332: data = 8'b00111100;	//   ****  
        12'h333: data = 8'b11000010;	// **    * 
        12'h334: data = 8'b00000010;	//       * 
        12'h335: data = 8'b00000000;	//         
        12'h336: data = 8'b00001100;	//     **  
        12'h337: data = 8'b00000010;	//       * 
        12'h338: data = 8'b11000010;	// **    * 
        12'h339: data = 8'b00111100;	//   ****  
        12'h33a: data = 8'b00000000;	//         
        12'h33b: data = 8'b00000000;	//         
        12'h33c: data = 8'b00000000;	//         
        12'h33d: data = 8'b00000000;	//         
        12'h33e: data = 8'b00000000;	//         
        12'h33f: data = 8'b00000000;	//         

    // code x34 (4)
        12'h340: data = 8'b00000000;	//         
        12'h341: data = 8'b00000000;	//         
        12'h342: data = 8'b00010000;	//    *    
        12'h343: data = 8'b00100000;	//   *     
        12'h344: data = 8'b11000000;	// **      
        12'h345: data = 8'b11000000;	// **      
        12'h346: data = 8'b11000100;	// **   *  
        12'h347: data = 8'b11000100;	// **   *  
        12'h348: data = 8'b11111110;	// ******* 
        12'h349: data = 8'b00000100;	//      *  
        12'h34a: data = 8'b00000000;	//         
        12'h34b: data = 8'b00000000;	//         
        12'h34c: data = 8'b00000000;	//         
        12'h34d: data = 8'b00000000;	//         
        12'h34e: data = 8'b00000000;	//         
        12'h34f: data = 8'b00000000;	//         

    // code x35 (5)
        12'h350: data = 8'b00000000;	//         
        12'h351: data = 8'b00000000;	//         
        12'h352: data = 8'b11111110;	// ******* 
        12'h353: data = 8'b11000000;	// **      
        12'h354: data = 8'b11000000;	// **      
        12'h355: data = 8'b01000000;	//  *      
        12'h356: data = 8'b00111100;	//   ****  
        12'h357: data = 8'b00000010;	//       * 
        12'h358: data = 8'b00000010;	//       * 
        12'h359: data = 8'b11111100;	// ******  
        12'h35a: data = 8'b00000000;	//         
        12'h35b: data = 8'b00000000;	//         
        12'h35c: data = 8'b00000000;	//         
        12'h35d: data = 8'b00000000;	//         
        12'h35e: data = 8'b00000000;	//         
        12'h35f: data = 8'b00000000;	//         

    // code x36 (6)
        12'h360: data = 8'b00000000;	//         
        12'h361: data = 8'b00000000;	//         
        12'h362: data = 8'b00111100;	//   ****  
        12'h363: data = 8'b00000010;	//       * 
        12'h364: data = 8'b11000000;	// **      
        12'h365: data = 8'b11000000;	// **      
        12'h366: data = 8'b11111100;	// ******  
        12'h367: data = 8'b11000010;	// **    * 
        12'h368: data = 8'b01000010;	//  *    * 
        12'h369: data = 8'b00111100;	//   ****  
        12'h36a: data = 8'b00000000;	//         
        12'h36b: data = 8'b00000000;	//         
        12'h36c: data = 8'b00000000;	//         
        12'h36d: data = 8'b00000000;	//         
        12'h36e: data = 8'b00000000;	//         
        12'h36f: data = 8'b00000000;	//         

    // code x37 (7)
        12'h370: data = 8'b00000000;	//         
        12'h371: data = 8'b00000000;	//         
        12'h372: data = 8'b11111100;	// ******  
        12'h373: data = 8'b00000010;	//       * 
        12'h374: data = 8'b00000010;	//       * 
        12'h375: data = 8'b00000010;	//       * 
        12'h376: data = 8'b00011110;	//    **** 
        12'h377: data = 8'b00000010;	//       * 
        12'h378: data = 8'b00000010;	//       * 
        12'h379: data = 8'b00000010;	//       * 
        12'h37a: data = 8'b00000000;	//         
        12'h37b: data = 8'b00000000;	//         
        12'h37c: data = 8'b00000000;	//         
        12'h37d: data = 8'b00000000;	//         
        12'h37e: data = 8'b00000000;	//         
        12'h37f: data = 8'b00000000;	//         

    // code x38 (8)
        12'h380: data = 8'b00000000;	//         
        12'h381: data = 8'b00000000;	//         
        12'h382: data = 8'b00111100;	//   ****  
        12'h383: data = 8'b11000010;	// **    * 
        12'h384: data = 8'b11000010;	// **    * 
        12'h385: data = 8'b00000000;	//         
        12'h386: data = 8'b00111100;	//   ****  
        12'h387: data = 8'b11000010;	// **    * 
        12'h388: data = 8'b11000010;	// **    * 
        12'h389: data = 8'b00111100;	//   ****  
        12'h38a: data = 8'b00000000;	//         
        12'h38b: data = 8'b00000000;	//         
        12'h38c: data = 8'b00000000;	//         
        12'h38d: data = 8'b00000000;	//         
        12'h38e: data = 8'b00000000;	//         
        12'h38f: data = 8'b00000000;	//         

    // code x39 (9)
        12'h390: data = 8'b00000000;	//         
        12'h391: data = 8'b00000000;	//         
        12'h392: data = 8'b00111100;	//   ****  
        12'h393: data = 8'b11000010;	// **    * 
        12'h394: data = 8'b11000010;	// **    * 
        12'h395: data = 8'b00000010;	//       * 
        12'h396: data = 8'b00111110;	//   ***** 
        12'h397: data = 8'b00000010;	//       * 
        12'h398: data = 8'b11000010;	// **    * 
        12'h399: data = 8'b00111100;	//   ****  
        12'h39a: data = 8'b00000000;	//         
        12'h39b: data = 8'b00000000;	//         
        12'h39c: data = 8'b00000000;	//         
        12'h39d: data = 8'b00000000;	//         
        12'h39e: data = 8'b00000000;	//         
        12'h39f: data = 8'b00000000;	//               

            default: data = 8'b00000000; // Default to zero
        endcase
 endmodule