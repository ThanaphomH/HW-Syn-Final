// *************************************************************
// Created by David J. Marion aka FPGA Dude
// A ROM containing patterns for ASCII values.
//
// Non-printable characters 00 - 1f, and 7f
// Printable characters 20 - 7e
//
// Not all character ROMs have been patterned.
// Only numbers, capital letters, some spec chars. 
//		Numbers       30 - 39
//   	Letters       41 - 5a 
//      (smiley face)   01
//		(space)         20
//		   .            2e
// 		   :            3a
//		   |	        7c	
//
// The 7-bit ASCII code for each character is used as
// the MSB of the address. The 4-bit LSB is the row value.
// *************************************************************

module ascii_rom(
        input clk, 
        input wire [10:0] addr,
        output reg [7:0] data
    );

    (* rom_style = "block" *) 

    reg [10:0] addr_reg;
    
    always @(posedge clk)
        addr_reg <= addr;
        
    always @*
        case(addr_reg)
    
    // code x41 (A)
        11'h410: data = 8'b00000000;	//         
        11'h411: data = 8'b00000000;	//         
        11'h412: data = 8'b00011000;	//    **   
        11'h413: data = 8'b00100100;	//   *  *  
        11'h414: data = 8'b11000010;	// **    * 
        11'h415: data = 8'b11000010;	// **    * 
        11'h416: data = 8'b11000010;	// **    * 
        11'h417: data = 8'b11111110;	// ******* 
        11'h418: data = 8'b11000010;	// **    * 
        11'h419: data = 8'b11000010;	// **    * 
        11'h41a: data = 8'b00000000;	//         
        11'h41b: data = 8'b00000000;	//         
        11'h41c: data = 8'b00000000;	//         
        11'h41d: data = 8'b00000000;	//         
        11'h41e: data = 8'b00000000;	//         
        11'h41f: data = 8'b00000000;	//         

    // code x42 (B)
        11'h420: data = 8'b00000000;	//         
        11'h421: data = 8'b00000000;	//         
        11'h422: data = 8'b11111100;	// ******  
        11'h423: data = 8'b11000010;	// **    * 
        11'h424: data = 8'b11000010;	// **    * 
        11'h425: data = 8'b11000000;	// **      
        11'h426: data = 8'b11111100;	// ******  
        11'h427: data = 8'b11000010;	// **    * 
        11'h428: data = 8'b11000010;	// **    * 
        11'h429: data = 8'b11111100;	// ******  
        11'h42a: data = 8'b00000000;	//         
        11'h42b: data = 8'b00000000;	//         
        11'h42c: data = 8'b00000000;	//         
        11'h42d: data = 8'b00000000;	//         
        11'h42e: data = 8'b00000000;	//         
        11'h42f: data = 8'b00000000;	//         

    // code x43 (C)
        11'h430: data = 8'b00000000;	//         
        11'h431: data = 8'b00000000;	//         
        11'h432: data = 8'b00111100;	//   ****  
        11'h433: data = 8'b00000010;	//       * 
        11'h434: data = 8'b11000010;	// **    * 
        11'h435: data = 8'b11000000;	// **      
        11'h436: data = 8'b11000000;	// **      
        11'h437: data = 8'b11000010;	// **    * 
        11'h438: data = 8'b11000010;	// **    * 
        11'h439: data = 8'b00111100;	//   ****  
        11'h43a: data = 8'b00000000;	//         
        11'h43b: data = 8'b00000000;	//         
        11'h43c: data = 8'b00000000;	//         
        11'h43d: data = 8'b00000000;	//         
        11'h43e: data = 8'b00000000;	//         
        11'h43f: data = 8'b00000000;	//         

    // code x44 (D)
        11'h440: data = 8'b00000000;	//         
        11'h441: data = 8'b00000000;	//         
        11'h442: data = 8'b11111000;	// *****   
        11'h443: data = 8'b11000100;	// **   *  
        11'h444: data = 8'b11000010;	// **    * 
        11'h445: data = 8'b11000010;	// **    * 
        11'h446: data = 8'b11000010;	// **    * 
        11'h447: data = 8'b11000010;	// **    * 
        11'h448: data = 8'b11000100;	// **   *  
        11'h449: data = 8'b11111000;	// *****   
        11'h44a: data = 8'b00000000;	//         
        11'h44b: data = 8'b00000000;	//         
        11'h44c: data = 8'b00000000;	//         
        11'h44d: data = 8'b00000000;	//         
        11'h44e: data = 8'b00000000;	//         
        11'h44f: data = 8'b00000000;	//         

    // code x45 (E)
        11'h450: data = 8'b00000000;	//         
        11'h451: data = 8'b00000000;	//         
        11'h452: data = 8'b11111100;	// ******  
        11'h453: data = 8'b11000000;	// **      
        11'h454: data = 8'b11000000;	// **      
        11'h455: data = 8'b11000000;	// **      
        11'h456: data = 8'b11111000;	// *****   
        11'h457: data = 8'b11000000;	// **      
        11'h458: data = 8'b11000000;	// **      
        11'h459: data = 8'b11111100;	// ******  
        11'h45a: data = 8'b00000000;	//         
        11'h45b: data = 8'b00000000;	//         
        11'h45c: data = 8'b00000000;	//         
        11'h45d: data = 8'b00000000;	//         
        11'h45e: data = 8'b00000000;	//         
        11'h45f: data = 8'b00000000;	//         

    // code x46 (F)
        11'h460: data = 8'b00000000;	//         
        11'h461: data = 8'b00000000;	//         
        11'h462: data = 8'b11111100;	// ******  
        11'h463: data = 8'b11000000;	// **      
        11'h464: data = 8'b11000000;	// **      
        11'h465: data = 8'b11000000;	// **      
        11'h466: data = 8'b11111000;	// *****   
        11'h467: data = 8'b11000000;	// **      
        11'h468: data = 8'b11000000;	// **      
        11'h469: data = 8'b11000000;	// **      
        11'h46a: data = 8'b00000000;	//         
        11'h46b: data = 8'b00000000;	//         
        11'h46c: data = 8'b00000000;	//         
        11'h46d: data = 8'b00000000;	//         
        11'h46e: data = 8'b00000000;	//         
        11'h46f: data = 8'b00000000;	//         

    // code x47 (G)
        11'h470: data = 8'b00000000;	//         
        11'h471: data = 8'b00000000;	//         
        11'h472: data = 8'b00111100;	//   ****  
        11'h473: data = 8'b00000010;	//       * 
        11'h474: data = 8'b11000000;	// **      
        11'h475: data = 8'b11000000;	// **      
        11'h476: data = 8'b11000110;	// **   ** 
        11'h477: data = 8'b11000010;	// **    * 
        11'h478: data = 8'b11000010;	// **    * 
        11'h479: data = 8'b00111100;	//   ****  
        11'h47a: data = 8'b00000000;	//         
        11'h47b: data = 8'b00000000;	//         
        11'h47c: data = 8'b00000000;	//         
        11'h47d: data = 8'b00000000;	//         
        11'h47e: data = 8'b00000000;	//         
        11'h47f: data = 8'b00000000;	//         

    // code x48 (H)
        11'h480: data = 8'b00000000;	//         
        11'h481: data = 8'b00000000;	//         
        11'h482: data = 8'b11000010;	// **    * 
        11'h483: data = 8'b11000010;	// **    * 
        11'h484: data = 8'b11000010;	// **    * 
        11'h485: data = 8'b11000010;	// **    * 
        11'h486: data = 8'b11111110;	// ******* 
        11'h487: data = 8'b11000010;	// **    * 
        11'h488: data = 8'b11000010;	// **    * 
        11'h489: data = 8'b11000010;	// **    * 
        11'h48a: data = 8'b00000000;	//         
        11'h48b: data = 8'b00000000;	//         
        11'h48c: data = 8'b00000000;	//         
        11'h48d: data = 8'b00000000;	//         
        11'h48e: data = 8'b00000000;	//         
        11'h48f: data = 8'b00000000;	//         

    // code x49 (I)
        11'h490: data = 8'b00000000;	//         
        11'h491: data = 8'b00000000;	//         
        11'h492: data = 8'b11000000;	// **      
        11'h493: data = 8'b11000000;	// **      
        11'h494: data = 8'b11000000;	// **      
        11'h495: data = 8'b11000000;	// **      
        11'h496: data = 8'b11000000;	// **      
        11'h497: data = 8'b11000000;	// **      
        11'h498: data = 8'b11000000;	// **      
        11'h499: data = 8'b11000000;	// **      
        11'h49a: data = 8'b00000000;	//         
        11'h49b: data = 8'b00000000;	//         
        11'h49c: data = 8'b00000000;	//         
        11'h49d: data = 8'b00000000;	//         
        11'h49e: data = 8'b00000000;	//         
        11'h49f: data = 8'b00000000;	//         

    // code x4a (J)
        11'h4a0: data = 8'b00000000;	//         
        11'h4a1: data = 8'b00000000;	//         
        11'h4a2: data = 8'b00010000;	//    *    
        11'h4a3: data = 8'b00010000;	//    *    
        11'h4a4: data = 8'b00010000;	//    *    
        11'h4a5: data = 8'b00010000;	//    *    
        11'h4a6: data = 8'b00010000;	//    *    
        11'h4a7: data = 8'b00010000;	//    *    
        11'h4a8: data = 8'b00010000;	//    *    
        11'h4a9: data = 8'b11100000;	// ***     
        11'h4aa: data = 8'b00000000;	//         
        11'h4ab: data = 8'b00000000;	//         
        11'h4ac: data = 8'b00000000;	//         
        11'h4ad: data = 8'b00000000;	//         
        11'h4ae: data = 8'b00000000;	//         
        11'h4af: data = 8'b00000000;	//         

    // code x4b (K)
        11'h4b0: data = 8'b00000000;	//         
        11'h4b1: data = 8'b00000000;	//         
        11'h4b2: data = 8'b11000010;	// **    * 
        11'h4b3: data = 8'b11000100;	// **   *  
        11'h4b4: data = 8'b11111000;	// *****   
        11'h4b5: data = 8'b11000100;	// **   *  
        11'h4b6: data = 8'b11000100;	// **   *  
        11'h4b7: data = 8'b11000010;	// **    * 
        11'h4b8: data = 8'b11000010;	// **    * 
        11'h4b9: data = 8'b11000010;	// **    * 
        11'h4ba: data = 8'b00000000;	//         
        11'h4bb: data = 8'b00000000;	//         
        11'h4bc: data = 8'b00000000;	//         
        11'h4bd: data = 8'b00000000;	//         
        11'h4be: data = 8'b00000000;	//         
        11'h4bf: data = 8'b00000000;	//         

    // code x4c (L)
        11'h4c0: data = 8'b00000000;	//         
        11'h4c1: data = 8'b00000000;	//         
        11'h4c2: data = 8'b11000000;	// **      
        11'h4c3: data = 8'b11000000;	// **      
        11'h4c4: data = 8'b11000000;	// **      
        11'h4c5: data = 8'b11000000;	// **      
        11'h4c6: data = 8'b11000000;	// **      
        11'h4c7: data = 8'b11000000;	// **      
        11'h4c8: data = 8'b11000000;	// **      
        11'h4c9: data = 8'b11111100;	// ******  
        11'h4ca: data = 8'b00000000;	//         
        11'h4cb: data = 8'b00000000;	//         
        11'h4cc: data = 8'b00000000;	//         
        11'h4cd: data = 8'b00000000;	//         
        11'h4ce: data = 8'b00000000;	//         
        11'h4cf: data = 8'b00000000;	//         

    // code x4d (M)
        11'h4d0: data = 8'b00000000;	//         
        11'h4d1: data = 8'b00000000;	//         
        11'h4d2: data = 8'b11100011;	// ***   **
        11'h4d3: data = 8'b11001001;	// **  *  *
        11'h4d4: data = 8'b11001001;	// **  *  *
        11'h4d5: data = 8'b11001001;	// **  *  *
        11'h4d6: data = 8'b11000001;	// **     *
        11'h4d7: data = 8'b11000001;	// **     *
        11'h4d8: data = 8'b11000001;	// **     *
        11'h4d9: data = 8'b11000001;	// **     *
        11'h4da: data = 8'b00000000;	//         
        11'h4db: data = 8'b00000000;	//         
        11'h4dc: data = 8'b00000000;	//         
        11'h4dd: data = 8'b00000000;	//         
        11'h4de: data = 8'b00000000;	//         
        11'h4df: data = 8'b00000000;	//         

    // code x4e (N)
        11'h4e0: data = 8'b00000000;	//         
        11'h4e1: data = 8'b00000000;	//         
        11'h4e2: data = 8'b11100010;	// ***   * 
        11'h4e3: data = 8'b11000010;	// **    * 
        11'h4e4: data = 8'b11000110;	// **   ** 
        11'h4e5: data = 8'b11000010;	// **    * 
        11'h4e6: data = 8'b11000010;	// **    * 
        11'h4e7: data = 8'b11000010;	// **    * 
        11'h4e8: data = 8'b11000010;	// **    * 
        11'h4e9: data = 8'b11000010;	// **    * 
        11'h4ea: data = 8'b00000000;	//         
        11'h4eb: data = 8'b00000000;	//         
        11'h4ec: data = 8'b00000000;	//         
        11'h4ed: data = 8'b00000000;	//         
        11'h4ee: data = 8'b00000000;	//         
        11'h4ef: data = 8'b00000000;	//         

    // code x4f (O)
        11'h4f0: data = 8'b00000000;	//         
        11'h4f1: data = 8'b00000000;	//         
        11'h4f2: data = 8'b00111100;	//   ****  
        11'h4f3: data = 8'b11000010;	// **    * 
        11'h4f4: data = 8'b11000010;	// **    * 
        11'h4f5: data = 8'b11000010;	// **    * 
        11'h4f6: data = 8'b11000010;	// **    * 
        11'h4f7: data = 8'b11000010;	// **    * 
        11'h4f8: data = 8'b11000010;	// **    * 
        11'h4f9: data = 8'b00111100;	//   ****  
        11'h4fa: data = 8'b00000000;	//         
        11'h4fb: data = 8'b00000000;	//         
        11'h4fc: data = 8'b00000000;	//         
        11'h4fd: data = 8'b00000000;	//         
        11'h4fe: data = 8'b00000000;	//         
        11'h4ff: data = 8'b00000000;	//         

    // code x50 (P)
        11'h500: data = 8'b00000000;	//         
        11'h501: data = 8'b00000000;	//         
        11'h502: data = 8'b11111100;	// ******  
        11'h503: data = 8'b11000010;	// **    * 
        11'h504: data = 8'b11000010;	// **    * 
        11'h505: data = 8'b11111100;	// ******  
        11'h506: data = 8'b11000000;	// **      
        11'h507: data = 8'b11000000;	// **      
        11'h508: data = 8'b11000000;	// **      
        11'h509: data = 8'b11000000;	// **      
        11'h50a: data = 8'b00000000;	//         
        11'h50b: data = 8'b00000000;	//         
        11'h50c: data = 8'b00000000;	//         
        11'h50d: data = 8'b00000000;	//         
        11'h50e: data = 8'b00000000;	//         
        11'h50f: data = 8'b00000000;	//         

    // code x51 (Q)
        11'h510: data = 8'b00000000;	//         
        11'h511: data = 8'b00000000;	//         
        11'h512: data = 8'b00111100;	//   ****  
        11'h513: data = 8'b11000010;	// **    * 
        11'h514: data = 8'b11000010;	// **    * 
        11'h515: data = 8'b11000010;	// **    * 
        11'h516: data = 8'b11000010;	// **    * 
        11'h517: data = 8'b11000010;	// **    * 
        11'h518: data = 8'b11000010;	// **    * 
        11'h519: data = 8'b00111100;	//   ****  
        11'h51a: data = 8'b00000000;	//         
        11'h51b: data = 8'b00000000;	//         
        11'h51c: data = 8'b00000000;	//         
        11'h51d: data = 8'b00000000;	//         
        11'h51e: data = 8'b00000000;	//         
        11'h51f: data = 8'b00000000;	//         

    // code x52 (R)
        11'h520: data = 8'b00000000;	//         
        11'h521: data = 8'b00000000;	//         
        11'h522: data = 8'b11111100;	// ******  
        11'h523: data = 8'b11000010;	// **    * 
        11'h524: data = 8'b11000010;	// **    * 
        11'h525: data = 8'b11000000;	// **      
        11'h526: data = 8'b11111100;	// ******  
        11'h527: data = 8'b11000010;	// **    * 
        11'h528: data = 8'b11000010;	// **    * 
        11'h529: data = 8'b11000010;	// **    * 
        11'h52a: data = 8'b00000000;	//         
        11'h52b: data = 8'b00000000;	//         
        11'h52c: data = 8'b00000000;	//         
        11'h52d: data = 8'b00000000;	//         
        11'h52e: data = 8'b00000000;	//         
        11'h52f: data = 8'b00000000;	//         

    // code x53 (S)
        11'h530: data = 8'b00000000;	//         
        11'h531: data = 8'b00000000;	//         
        11'h532: data = 8'b00111100;	//   ****  
        11'h533: data = 8'b11000010;	// **    * 
        11'h534: data = 8'b11000000;	// **      
        11'h535: data = 8'b00000000;	//         
        11'h536: data = 8'b00111100;	//   ****  
        11'h537: data = 8'b00000010;	//       * 
        11'h538: data = 8'b11000010;	// **    * 
        11'h539: data = 8'b00111100;	//   ****  
        11'h53a: data = 8'b00000000;	//         
        11'h53b: data = 8'b00000000;	//         
        11'h53c: data = 8'b00000000;	//         
        11'h53d: data = 8'b00000000;	//         
        11'h53e: data = 8'b00000000;	//         
        11'h53f: data = 8'b00000000;	//         

    // code x54 (T)
        11'h540: data = 8'b00000000;	//         
        11'h541: data = 8'b00000000;	//         
        11'h542: data = 8'b11111100;	// ******  
        11'h543: data = 8'b00010000;	//    *    
        11'h544: data = 8'b00010000;	//    *    
        11'h545: data = 8'b00010000;	//    *    
        11'h546: data = 8'b00010000;	//    *    
        11'h547: data = 8'b00010000;	//    *    
        11'h548: data = 8'b00010000;	//    *    
        11'h549: data = 8'b00010000;	//    *    
        11'h54a: data = 8'b00000000;	//         
        11'h54b: data = 8'b00000000;	//         
        11'h54c: data = 8'b00000000;	//         
        11'h54d: data = 8'b00000000;	//         
        11'h54e: data = 8'b00000000;	//         
        11'h54f: data = 8'b00000000;	//         

    // code x55 (U)
        11'h550: data = 8'b00000000;	//         
        11'h551: data = 8'b00000000;	//         
        11'h552: data = 8'b11000010;	// **    * 
        11'h553: data = 8'b11000010;	// **    * 
        11'h554: data = 8'b11000010;	// **    * 
        11'h555: data = 8'b11000010;	// **    * 
        11'h556: data = 8'b11000010;	// **    * 
        11'h557: data = 8'b11000010;	// **    * 
        11'h558: data = 8'b11000010;	// **    * 
        11'h559: data = 8'b00111100;	//   ****  
        11'h55a: data = 8'b00000000;	//         
        11'h55b: data = 8'b00000000;	//         
        11'h55c: data = 8'b00000000;	//         
        11'h55d: data = 8'b00000000;	//         
        11'h55e: data = 8'b00000000;	//         
        11'h55f: data = 8'b00000000;	//         

    // code x56 (V)
        11'h560: data = 8'b00000000;	//         
        11'h561: data = 8'b00000000;	//         
        11'h562: data = 8'b11000010;	// **    * 
        11'h563: data = 8'b11000010;	// **    * 
        11'h564: data = 8'b11000010;	// **    * 
        11'h565: data = 8'b11000010;	// **    * 
        11'h566: data = 8'b11000010;	// **    * 
        11'h567: data = 8'b11000010;	// **    * 
        11'h568: data = 8'b00100100;	//   *  *  
        11'h569: data = 8'b00011000;	//    **   
        11'h56a: data = 8'b00000000;	//         
        11'h56b: data = 8'b00000000;	//         
        11'h56c: data = 8'b00000000;	//         
        11'h56d: data = 8'b00000000;	//         
        11'h56e: data = 8'b00000000;	//         
        11'h56f: data = 8'b00000000;	//         

    // code x57 (W)
        11'h570: data = 8'b00000000;	//         
        11'h571: data = 8'b00000000;	//         
        11'h572: data = 8'b11000001;	// **     *
        11'h573: data = 8'b11000001;	// **     *
        11'h574: data = 8'b11000001;	// **     *
        11'h575: data = 8'b11001001;	// **  *  *
        11'h576: data = 8'b11001001;	// **  *  *
        11'h577: data = 8'b11001001;	// **  *  *
        11'h578: data = 8'b11001001;	// **  *  *
        11'h579: data = 8'b00100010;	//   *   * 
        11'h57a: data = 8'b00000000;	//         
        11'h57b: data = 8'b00000000;	//         
        11'h57c: data = 8'b00000000;	//         
        11'h57d: data = 8'b00000000;	//         
        11'h57e: data = 8'b00000000;	//         
        11'h57f: data = 8'b00000000;	//         

    // code x58 (X)
        11'h580: data = 8'b00000000;	//         
        11'h581: data = 8'b00000000;	//         
        11'h582: data = 8'b00000100;	//      *  
        11'h583: data = 8'b11000100;	// **   *  
        11'h584: data = 8'b00000000;	//         
        11'h585: data = 8'b00010000;	//    *    
        11'h586: data = 8'b00010000;	//    *    
        11'h587: data = 8'b00000000;	//         
        11'h588: data = 8'b11000100;	// **   *  
        11'h589: data = 8'b11000100;	// **   *  
        11'h58a: data = 8'b00000000;	//         
        11'h58b: data = 8'b00000000;	//         
        11'h58c: data = 8'b00000000;	//         
        11'h58d: data = 8'b00000000;	//         
        11'h58e: data = 8'b00000000;	//         
        11'h58f: data = 8'b00000000;	//         

    // code x59 (Y)
        11'h590: data = 8'b00000000;	//         
        11'h591: data = 8'b00000000;	//         
        11'h592: data = 8'b11000100;	// **   *  
        11'h593: data = 8'b11000100;	// **   *  
        11'h594: data = 8'b11000100;	// **   *  
        11'h595: data = 8'b00111000;	//   ***   
        11'h596: data = 8'b00010000;	//    *    
        11'h597: data = 8'b00010000;	//    *    
        11'h598: data = 8'b00010000;	//    *    
        11'h599: data = 8'b00010000;	//    *    
        11'h59a: data = 8'b00000000;	//         
        11'h59b: data = 8'b00000000;	//         
        11'h59c: data = 8'b00000000;	//         
        11'h59d: data = 8'b00000000;	//         
        11'h59e: data = 8'b00000000;	//         
        11'h59f: data = 8'b00000000;	//         

    // code x5a (Z)
        11'h5a0: data = 8'b00000000;	//         
        11'h5a1: data = 8'b00000000;	//         
        11'h5a2: data = 8'b11111100;	// ******  
        11'h5a3: data = 8'b00000100;	//      *  
        11'h5a4: data = 8'b00001000;	//     *   
        11'h5a5: data = 8'b00001000;	//     *   
        11'h5a6: data = 8'b00010000;	//    *    
        11'h5a7: data = 8'b00100000;	//   *     
        11'h5a8: data = 8'b11000000;	// **      
        11'h5a9: data = 8'b11111100;	// ******  
        11'h5aa: data = 8'b00000000;	//         
        11'h5ab: data = 8'b00000000;	//         
        11'h5ac: data = 8'b00000000;	//         
        11'h5ad: data = 8'b00000000;	//         
        11'h5ae: data = 8'b00000000;	//         
        11'h5af: data = 8'b00000000;	//         

    // code x61 (a)
        11'h610: data = 8'b00000000;	//         
        11'h611: data = 8'b00000000;	//         
        11'h612: data = 8'b00000000;	//         
        11'h613: data = 8'b00111100;	//   ****  
        11'h614: data = 8'b00000010;	//       * 
        11'h615: data = 8'b00000010;	//       * 
        11'h616: data = 8'b00111110;	//   ***** 
        11'h617: data = 8'b11000010;	// **    * 
        11'h618: data = 8'b11000010;	// **    * 
        11'h619: data = 8'b00111110;	//   ***** 
        11'h61a: data = 8'b00000000;	//         
        11'h61b: data = 8'b00000000;	//         
        11'h61c: data = 8'b00000000;	//         
        11'h61d: data = 8'b00000000;	//         
        11'h61e: data = 8'b00000000;	//         
        11'h61f: data = 8'b00000000;	//         

    // code x62 (b)
        11'h620: data = 8'b00000000;	//         
        11'h621: data = 8'b11000000;	// **      
        11'h622: data = 8'b11000000;	// **      
        11'h623: data = 8'b11111100;	// ******  
        11'h624: data = 8'b11000010;	// **    * 
        11'h625: data = 8'b11000010;	// **    * 
        11'h626: data = 8'b11000010;	// **    * 
        11'h627: data = 8'b11000010;	// **    * 
        11'h628: data = 8'b11000010;	// **    * 
        11'h629: data = 8'b11111100;	// ******  
        11'h62a: data = 8'b00000000;	//         
        11'h62b: data = 8'b00000000;	//         
        11'h62c: data = 8'b00000000;	//         
        11'h62d: data = 8'b00000000;	//         
        11'h62e: data = 8'b00000000;	//         
        11'h62f: data = 8'b00000000;	//         

    // code x63 (c)
        11'h630: data = 8'b00000000;	//         
        11'h631: data = 8'b00000000;	//         
        11'h632: data = 8'b00000000;	//         
        11'h633: data = 8'b00111100;	//   ****  
        11'h634: data = 8'b11000000;	// **      
        11'h635: data = 8'b11000010;	// **    * 
        11'h636: data = 8'b11000000;	// **      
        11'h637: data = 8'b11000000;	// **      
        11'h638: data = 8'b11000010;	// **    * 
        11'h639: data = 8'b00111100;	//   ****  
        11'h63a: data = 8'b00000000;	//         
        11'h63b: data = 8'b00000000;	//         
        11'h63c: data = 8'b00000000;	//         
        11'h63d: data = 8'b00000000;	//         
        11'h63e: data = 8'b00000000;	//         
        11'h63f: data = 8'b00000000;	//         

    // code x64 (d)
        11'h640: data = 8'b00000000;	//         
        11'h641: data = 8'b00000010;	//       * 
        11'h642: data = 8'b00000010;	//       * 
        11'h643: data = 8'b00111110;	//   ***** 
        11'h644: data = 8'b11000010;	// **    * 
        11'h645: data = 8'b11000010;	// **    * 
        11'h646: data = 8'b11000010;	// **    * 
        11'h647: data = 8'b11000010;	// **    * 
        11'h648: data = 8'b11000010;	// **    * 
        11'h649: data = 8'b00111110;	//   ***** 
        11'h64a: data = 8'b00000000;	//         
        11'h64b: data = 8'b00000000;	//         
        11'h64c: data = 8'b00000000;	//         
        11'h64d: data = 8'b00000000;	//         
        11'h64e: data = 8'b00000000;	//         
        11'h64f: data = 8'b00000000;	//         

    // code x65 (e)
        11'h650: data = 8'b00000000;	//         
        11'h651: data = 8'b00000000;	//         
        11'h652: data = 8'b00000000;	//         
        11'h653: data = 8'b00111100;	//   ****  
        11'h654: data = 8'b11000000;	// **      
        11'h655: data = 8'b11000010;	// **    * 
        11'h656: data = 8'b11000010;	// **    * 
        11'h657: data = 8'b11111100;	// ******  
        11'h658: data = 8'b11000000;	// **      
        11'h659: data = 8'b00111100;	//   ****  
        11'h65a: data = 8'b00000000;	//         
        11'h65b: data = 8'b00000000;	//         
        11'h65c: data = 8'b00000000;	//         
        11'h65d: data = 8'b00000000;	//         
        11'h65e: data = 8'b00000000;	//         
        11'h65f: data = 8'b00000000;	//         

    // code x66 (f)
        11'h660: data = 8'b00000000;	//         
        11'h661: data = 8'b00110000;	//   **    
        11'h662: data = 8'b11000000;	// **      
        11'h663: data = 8'b11000000;	// **      
        11'h664: data = 8'b11000000;	// **      
        11'h665: data = 8'b11110000;	// ****    
        11'h666: data = 8'b11000000;	// **      
        11'h667: data = 8'b11000000;	// **      
        11'h668: data = 8'b11000000;	// **      
        11'h669: data = 8'b11000000;	// **      
        11'h66a: data = 8'b00000000;	//         
        11'h66b: data = 8'b00000000;	//         
        11'h66c: data = 8'b00000000;	//         
        11'h66d: data = 8'b00000000;	//         
        11'h66e: data = 8'b00000000;	//         
        11'h66f: data = 8'b00000000;	//         

    // code x67 (g)
        11'h670: data = 8'b00000000;	//         
        11'h671: data = 8'b00000000;	//         
        11'h672: data = 8'b00000100;	//      *  
        11'h673: data = 8'b00111110;	//   ***** 
        11'h674: data = 8'b11000010;	// **    * 
        11'h675: data = 8'b11000010;	// **    * 
        11'h676: data = 8'b00000000;	//         
        11'h677: data = 8'b00111100;	//   ****  
        11'h678: data = 8'b00001000;	//     *   
        11'h679: data = 8'b00111100;	//   ****  
        11'h67a: data = 8'b11000010;	// **    * 
        11'h67b: data = 8'b11000010;	// **    * 
        11'h67c: data = 8'b00000000;	//         
        11'h67d: data = 8'b00000000;	//         
        11'h67e: data = 8'b00000000;	//         
        11'h67f: data = 8'b00000000;	//         

    // code x68 (h)
        11'h680: data = 8'b00000000;	//         
        11'h681: data = 8'b11000000;	// **      
        11'h682: data = 8'b11000000;	// **      
        11'h683: data = 8'b11111100;	// ******  
        11'h684: data = 8'b11000010;	// **    * 
        11'h685: data = 8'b11000010;	// **    * 
        11'h686: data = 8'b11000010;	// **    * 
        11'h687: data = 8'b11000010;	// **    * 
        11'h688: data = 8'b11000010;	// **    * 
        11'h689: data = 8'b11000010;	// **    * 
        11'h68a: data = 8'b00000000;	//         
        11'h68b: data = 8'b00000000;	//         
        11'h68c: data = 8'b00000000;	//         
        11'h68d: data = 8'b00000000;	//         
        11'h68e: data = 8'b00000000;	//         
        11'h68f: data = 8'b00000000;	//         

    // code x69 (i)
        11'h690: data = 8'b00000000;	//         
        11'h691: data = 8'b11000000;	// **      
        11'h692: data = 8'b00000000;	//         
        11'h693: data = 8'b00000000;	//         
        11'h694: data = 8'b11000000;	// **      
        11'h695: data = 8'b11000000;	// **      
        11'h696: data = 8'b11000000;	// **      
        11'h697: data = 8'b11000000;	// **      
        11'h698: data = 8'b11000000;	// **      
        11'h699: data = 8'b11000000;	// **      
        11'h69a: data = 8'b00000000;	//         
        11'h69b: data = 8'b00000000;	//         
        11'h69c: data = 8'b00000000;	//         
        11'h69d: data = 8'b00000000;	//         
        11'h69e: data = 8'b00000000;	//         
        11'h69f: data = 8'b00000000;	//         

    // code x6a (j)
        11'h6a0: data = 8'b00000000;	//         
        11'h6a1: data = 8'b11000000;	// **      
        11'h6a2: data = 8'b00000000;	//         
        11'h6a3: data = 8'b00000000;	//         
        11'h6a4: data = 8'b11000000;	// **      
        11'h6a5: data = 8'b11000000;	// **      
        11'h6a6: data = 8'b11000000;	// **      
        11'h6a7: data = 8'b11000000;	// **      
        11'h6a8: data = 8'b11000000;	// **      
        11'h6a9: data = 8'b11000000;	// **      
        11'h6aa: data = 8'b11000000;	// **      
        11'h6ab: data = 8'b10000000;	// *       
        11'h6ac: data = 8'b00000000;	//         
        11'h6ad: data = 8'b00000000;	//         
        11'h6ae: data = 8'b00000000;	//         
        11'h6af: data = 8'b00000000;	//         

    // code x6b (k)
        11'h6b0: data = 8'b00000000;	//         
        11'h6b1: data = 8'b11000000;	// **      
        11'h6b2: data = 8'b11000000;	// **      
        11'h6b3: data = 8'b11000100;	// **   *  
        11'h6b4: data = 8'b11001000;	// **  *   
        11'h6b5: data = 8'b11000000;	// **      
        11'h6b6: data = 8'b11110000;	// ****    
        11'h6b7: data = 8'b11001000;	// **  *   
        11'h6b8: data = 8'b11000100;	// **   *  
        11'h6b9: data = 8'b11000100;	// **   *  
        11'h6ba: data = 8'b00000000;	//         
        11'h6bb: data = 8'b00000000;	//         
        11'h6bc: data = 8'b00000000;	//         
        11'h6bd: data = 8'b00000000;	//         
        11'h6be: data = 8'b00000000;	//         
        11'h6bf: data = 8'b00000000;	//         

    // code x6c (l)
        11'h6c0: data = 8'b00000000;	//         
        11'h6c1: data = 8'b11000000;	// **      
        11'h6c2: data = 8'b11000000;	// **      
        11'h6c3: data = 8'b11000000;	// **      
        11'h6c4: data = 8'b11000000;	// **      
        11'h6c5: data = 8'b11000000;	// **      
        11'h6c6: data = 8'b11000000;	// **      
        11'h6c7: data = 8'b11000000;	// **      
        11'h6c8: data = 8'b11000000;	// **      
        11'h6c9: data = 8'b11000000;	// **      
        11'h6ca: data = 8'b00000000;	//         
        11'h6cb: data = 8'b00000000;	//         
        11'h6cc: data = 8'b00000000;	//         
        11'h6cd: data = 8'b00000000;	//         
        11'h6ce: data = 8'b00000000;	//         
        11'h6cf: data = 8'b00000000;	//         

    // code x6d (m)
        11'h6d0: data = 8'b00000000;	//         
        11'h6d1: data = 8'b00000000;	//         
        11'h6d2: data = 8'b00000000;	//         
        11'h6d3: data = 8'b11100010;	// ***   * 
        11'h6d4: data = 8'b11001001;	// **  *  *
        11'h6d5: data = 8'b11001001;	// **  *  *
        11'h6d6: data = 8'b11001001;	// **  *  *
        11'h6d7: data = 8'b11001001;	// **  *  *
        11'h6d8: data = 8'b11001001;	// **  *  *
        11'h6d9: data = 8'b11001001;	// **  *  *
        11'h6da: data = 8'b00000000;	//         
        11'h6db: data = 8'b00000000;	//         
        11'h6dc: data = 8'b00000000;	//         
        11'h6dd: data = 8'b00000000;	//         
        11'h6de: data = 8'b00000000;	//         
        11'h6df: data = 8'b00000000;	//         

    // code x6e (n)
        11'h6e0: data = 8'b00000000;	//         
        11'h6e1: data = 8'b00000000;	//         
        11'h6e2: data = 8'b00000000;	//         
        11'h6e3: data = 8'b11111100;	// ******  
        11'h6e4: data = 8'b11000010;	// **    * 
        11'h6e5: data = 8'b11000010;	// **    * 
        11'h6e6: data = 8'b11000010;	// **    * 
        11'h6e7: data = 8'b11000010;	// **    * 
        11'h6e8: data = 8'b11000010;	// **    * 
        11'h6e9: data = 8'b11000010;	// **    * 
        11'h6ea: data = 8'b00000000;	//         
        11'h6eb: data = 8'b00000000;	//         
        11'h6ec: data = 8'b00000000;	//         
        11'h6ed: data = 8'b00000000;	//         
        11'h6ee: data = 8'b00000000;	//         
        11'h6ef: data = 8'b00000000;	//         

    // code x6f (o)
        11'h6f0: data = 8'b00000000;	//         
        11'h6f1: data = 8'b00000000;	//         
        11'h6f2: data = 8'b00000000;	//         
        11'h6f3: data = 8'b00111100;	//   ****  
        11'h6f4: data = 8'b11000010;	// **    * 
        11'h6f5: data = 8'b11000010;	// **    * 
        11'h6f6: data = 8'b11000010;	// **    * 
        11'h6f7: data = 8'b11000010;	// **    * 
        11'h6f8: data = 8'b11000010;	// **    * 
        11'h6f9: data = 8'b00111100;	//   ****  
        11'h6fa: data = 8'b00000000;	//         
        11'h6fb: data = 8'b00000000;	//         
        11'h6fc: data = 8'b00000000;	//         
        11'h6fd: data = 8'b00000000;	//         
        11'h6fe: data = 8'b00000000;	//         
        11'h6ff: data = 8'b00000000;	//         

    // code x70 (p)
        11'h700: data = 8'b00000000;	//         
        11'h701: data = 8'b00000000;	//         
        11'h702: data = 8'b00000000;	//         
        11'h703: data = 8'b11111100;	// ******  
        11'h704: data = 8'b11000010;	// **    * 
        11'h705: data = 8'b11000010;	// **    * 
        11'h706: data = 8'b11000010;	// **    * 
        11'h707: data = 8'b11000010;	// **    * 
        11'h708: data = 8'b11000010;	// **    * 
        11'h709: data = 8'b11111100;	// ******  
        11'h70a: data = 8'b11000000;	// **      
        11'h70b: data = 8'b11000000;	// **      
        11'h70c: data = 8'b00000000;	//         
        11'h70d: data = 8'b00000000;	//         
        11'h70e: data = 8'b00000000;	//         
        11'h70f: data = 8'b00000000;	//         

    // code x71 (q)
        11'h710: data = 8'b00000000;	//         
        11'h711: data = 8'b00000000;	//         
        11'h712: data = 8'b00000000;	//         
        11'h713: data = 8'b00111110;	//   ***** 
        11'h714: data = 8'b11000010;	// **    * 
        11'h715: data = 8'b11000010;	// **    * 
        11'h716: data = 8'b11000010;	// **    * 
        11'h717: data = 8'b11000010;	// **    * 
        11'h718: data = 8'b11000010;	// **    * 
        11'h719: data = 8'b00111110;	//   ***** 
        11'h71a: data = 8'b00000010;	//       * 
        11'h71b: data = 8'b00000010;	//       * 
        11'h71c: data = 8'b00000000;	//         
        11'h71d: data = 8'b00000000;	//         
        11'h71e: data = 8'b00000000;	//         
        11'h71f: data = 8'b00000000;	//         

    // code x72 (r)
        11'h720: data = 8'b00000000;	//         
        11'h721: data = 8'b00000000;	//         
        11'h722: data = 8'b00000000;	//         
        11'h723: data = 8'b11111000;	// *****   
        11'h724: data = 8'b11000100;	// **   *  
        11'h725: data = 8'b11000000;	// **      
        11'h726: data = 8'b11000000;	// **      
        11'h727: data = 8'b11000000;	// **      
        11'h728: data = 8'b11000000;	// **      
        11'h729: data = 8'b11000000;	// **      
        11'h72a: data = 8'b00000000;	//         
        11'h72b: data = 8'b00000000;	//         
        11'h72c: data = 8'b00000000;	//         
        11'h72d: data = 8'b00000000;	//         
        11'h72e: data = 8'b00000000;	//         
        11'h72f: data = 8'b00000000;	//         

    // code x73 (s)
        11'h730: data = 8'b00000000;	//         
        11'h731: data = 8'b00000000;	//         
        11'h732: data = 8'b00000000;	//         
        11'h733: data = 8'b00111100;	//   ****  
        11'h734: data = 8'b11000000;	// **      
        11'h735: data = 8'b00000000;	//         
        11'h736: data = 8'b00111000;	//   ***   
        11'h737: data = 8'b00000100;	//      *  
        11'h738: data = 8'b00000100;	//      *  
        11'h739: data = 8'b11111000;	// *****   
        11'h73a: data = 8'b00000000;	//         
        11'h73b: data = 8'b00000000;	//         
        11'h73c: data = 8'b00000000;	//         
        11'h73d: data = 8'b00000000;	//         
        11'h73e: data = 8'b00000000;	//         
        11'h73f: data = 8'b00000000;	//         

    // code x74 (t)
        11'h740: data = 8'b00000000;	//         
        11'h741: data = 8'b00100000;	//   *     
        11'h742: data = 8'b00100000;	//   *     
        11'h743: data = 8'b11110000;	// ****    
        11'h744: data = 8'b00100000;	//   *     
        11'h745: data = 8'b00100000;	//   *     
        11'h746: data = 8'b00100000;	//   *     
        11'h747: data = 8'b00100000;	//   *     
        11'h748: data = 8'b00100000;	//   *     
        11'h749: data = 8'b00010000;	//    *    
        11'h74a: data = 8'b00000000;	//         
        11'h74b: data = 8'b00000000;	//         
        11'h74c: data = 8'b00000000;	//         
        11'h74d: data = 8'b00000000;	//         
        11'h74e: data = 8'b00000000;	//         
        11'h74f: data = 8'b00000000;	//         

    // code x75 (u)
        11'h750: data = 8'b00000000;	//         
        11'h751: data = 8'b00000000;	//         
        11'h752: data = 8'b00000000;	//         
        11'h753: data = 8'b11000010;	// **    * 
        11'h754: data = 8'b11000010;	// **    * 
        11'h755: data = 8'b11000010;	// **    * 
        11'h756: data = 8'b11000010;	// **    * 
        11'h757: data = 8'b11000010;	// **    * 
        11'h758: data = 8'b11000010;	// **    * 
        11'h759: data = 8'b00111110;	//   ***** 
        11'h75a: data = 8'b00000000;	//         
        11'h75b: data = 8'b00000000;	//         
        11'h75c: data = 8'b00000000;	//         
        11'h75d: data = 8'b00000000;	//         
        11'h75e: data = 8'b00000000;	//         
        11'h75f: data = 8'b00000000;	//         

    // code x76 (v)
        11'h760: data = 8'b00000000;	//         
        11'h761: data = 8'b00000000;	//         
        11'h762: data = 8'b00000000;	//         
        11'h763: data = 8'b11000010;	// **    * 
        11'h764: data = 8'b11000010;	// **    * 
        11'h765: data = 8'b11000010;	// **    * 
        11'h766: data = 8'b11000010;	// **    * 
        11'h767: data = 8'b11000010;	// **    * 
        11'h768: data = 8'b00100100;	//   *  *  
        11'h769: data = 8'b00011000;	//    **   
        11'h76a: data = 8'b00000000;	//         
        11'h76b: data = 8'b00000000;	//         
        11'h76c: data = 8'b00000000;	//         
        11'h76d: data = 8'b00000000;	//         
        11'h76e: data = 8'b00000000;	//         
        11'h76f: data = 8'b00000000;	//         

    // code x77 (w)
        11'h770: data = 8'b00000000;	//         
        11'h771: data = 8'b00000000;	//         
        11'h772: data = 8'b00000000;	//         
        11'h773: data = 8'b11000010;	// **    * 
        11'h774: data = 8'b11000010;	// **    * 
        11'h775: data = 8'b11000010;	// **    * 
        11'h776: data = 8'b11000010;	// **    * 
        11'h777: data = 8'b11000010;	// **    * 
        11'h778: data = 8'b11000010;	// **    * 
        11'h779: data = 8'b00100100;	//   *  *  
        11'h77a: data = 8'b00000000;	//         
        11'h77b: data = 8'b00000000;	//         
        11'h77c: data = 8'b00000000;	//         
        11'h77d: data = 8'b00000000;	//         
        11'h77e: data = 8'b00000000;	//         
        11'h77f: data = 8'b00000000;	//         

    // code x78 (x)
        11'h780: data = 8'b00000000;	//         
        11'h781: data = 8'b00000000;	//         
        11'h782: data = 8'b00000000;	//         
        11'h783: data = 8'b11000000;	// **      
        11'h784: data = 8'b00100100;	//   *  *  
        11'h785: data = 8'b00000000;	//         
        11'h786: data = 8'b00011000;	//    **   
        11'h787: data = 8'b00100100;	//   *  *  
        11'h788: data = 8'b11000010;	// **    * 
        11'h789: data = 8'b11000010;	// **    * 
        11'h78a: data = 8'b00000000;	//         
        11'h78b: data = 8'b00000000;	//         
        11'h78c: data = 8'b00000000;	//         
        11'h78d: data = 8'b00000000;	//         
        11'h78e: data = 8'b00000000;	//         
        11'h78f: data = 8'b00000000;	//         

    // code x79 (y)
        11'h790: data = 8'b00000000;	//         
        11'h791: data = 8'b00000000;	//         
        11'h792: data = 8'b00000000;	//         
        11'h793: data = 8'b11000010;	// **    * 
        11'h794: data = 8'b11000010;	// **    * 
        11'h795: data = 8'b11000010;	// **    * 
        11'h796: data = 8'b11000010;	// **    * 
        11'h797: data = 8'b11000010;	// **    * 
        11'h798: data = 8'b11000010;	// **    * 
        11'h799: data = 8'b00111110;	//   ***** 
        11'h79a: data = 8'b00000010;	//       * 
        11'h79b: data = 8'b00111100;	//   ****  
        11'h79c: data = 8'b00000000;	//         
        11'h79d: data = 8'b00000000;	//         
        11'h79e: data = 8'b00000000;	//         
        11'h79f: data = 8'b00000000;	//         

    // code x7a (z)
        11'h7a0: data = 8'b00000000;	//         
        11'h7a1: data = 8'b00000000;	//         
        11'h7a2: data = 8'b00000000;	//         
        11'h7a3: data = 8'b00000000;	//         
        11'h7a4: data = 8'b00001000;	//     *   
        11'h7a5: data = 8'b00010000;	//    *    
        11'h7a6: data = 8'b00010000;	//    *    
        11'h7a7: data = 8'b01000000;	//  *      
        11'h7a8: data = 8'b11000000;	// **      
        11'h7a9: data = 8'b11111000;	// *****   
        11'h7aa: data = 8'b00000000;	//         
        11'h7ab: data = 8'b00000000;	//         
        11'h7ac: data = 8'b00000000;	//         
        11'h7ad: data = 8'b00000000;	//         
        11'h7ae: data = 8'b00000000;	//         
        11'h7af: data = 8'b00000000;	//         

    // code x30 (0)
        11'h300: data = 8'b00000000;	//         
        11'h301: data = 8'b00000000;	//         
        11'h302: data = 8'b00111100;	//   ****  
        11'h303: data = 8'b11000010;	// **    * 
        11'h304: data = 8'b11000010;	// **    * 
        11'h305: data = 8'b11000010;	// **    * 
        11'h306: data = 8'b11000110;	// **   ** 
        11'h307: data = 8'b11000010;	// **    * 
        11'h308: data = 8'b11100010;	// ***   * 
        11'h309: data = 8'b00111100;	//   ****  
        11'h30a: data = 8'b00000000;	//         
        11'h30b: data = 8'b00000000;	//         
        11'h30c: data = 8'b00000000;	//         
        11'h30d: data = 8'b00000000;	//         
        11'h30e: data = 8'b00000000;	//         
        11'h30f: data = 8'b00000000;	//         

    // code x31 (1)
        11'h310: data = 8'b00000000;	//         
        11'h311: data = 8'b00000000;	//         
        11'h312: data = 8'b00100000;	//   *     
        11'h313: data = 8'b11100000;	// ***     
        11'h314: data = 8'b00100000;	//   *     
        11'h315: data = 8'b00100000;	//   *     
        11'h316: data = 8'b00100000;	//   *     
        11'h317: data = 8'b00100000;	//   *     
        11'h318: data = 8'b00100000;	//   *     
        11'h319: data = 8'b11110000;	// ****    
        11'h31a: data = 8'b00000000;	//         
        11'h31b: data = 8'b00000000;	//         
        11'h31c: data = 8'b00000000;	//         
        11'h31d: data = 8'b00000000;	//         
        11'h31e: data = 8'b00000000;	//         
        11'h31f: data = 8'b00000000;	//         

    // code x32 (2)
        11'h320: data = 8'b00000000;	//         
        11'h321: data = 8'b00000000;	//         
        11'h322: data = 8'b00111100;	//   ****  
        11'h323: data = 8'b11000010;	// **    * 
        11'h324: data = 8'b00000010;	//       * 
        11'h325: data = 8'b00000010;	//       * 
        11'h326: data = 8'b00011100;	//    ***  
        11'h327: data = 8'b00100000;	//   *     
        11'h328: data = 8'b11000000;	// **      
        11'h329: data = 8'b11111110;	// ******* 
        11'h32a: data = 8'b00000000;	//         
        11'h32b: data = 8'b00000000;	//         
        11'h32c: data = 8'b00000000;	//         
        11'h32d: data = 8'b00000000;	//         
        11'h32e: data = 8'b00000000;	//         
        11'h32f: data = 8'b00000000;	//         

    // code x33 (3)
        11'h330: data = 8'b00000000;	//         
        11'h331: data = 8'b00000000;	//         
        11'h332: data = 8'b00111100;	//   ****  
        11'h333: data = 8'b11000010;	// **    * 
        11'h334: data = 8'b00000010;	//       * 
        11'h335: data = 8'b00000000;	//         
        11'h336: data = 8'b00001100;	//     **  
        11'h337: data = 8'b00000010;	//       * 
        11'h338: data = 8'b11000010;	// **    * 
        11'h339: data = 8'b00111100;	//   ****  
        11'h33a: data = 8'b00000000;	//         
        11'h33b: data = 8'b00000000;	//         
        11'h33c: data = 8'b00000000;	//         
        11'h33d: data = 8'b00000000;	//         
        11'h33e: data = 8'b00000000;	//         
        11'h33f: data = 8'b00000000;	//         

    // code x34 (4)
        11'h340: data = 8'b00000000;	//         
        11'h341: data = 8'b00000000;	//         
        11'h342: data = 8'b00010000;	//    *    
        11'h343: data = 8'b00100000;	//   *     
        11'h344: data = 8'b11000000;	// **      
        11'h345: data = 8'b11000000;	// **      
        11'h346: data = 8'b11000100;	// **   *  
        11'h347: data = 8'b11000100;	// **   *  
        11'h348: data = 8'b11111110;	// ******* 
        11'h349: data = 8'b00000100;	//      *  
        11'h34a: data = 8'b00000000;	//         
        11'h34b: data = 8'b00000000;	//         
        11'h34c: data = 8'b00000000;	//         
        11'h34d: data = 8'b00000000;	//         
        11'h34e: data = 8'b00000000;	//         
        11'h34f: data = 8'b00000000;	//         

    // code x35 (5)
        11'h350: data = 8'b00000000;	//         
        11'h351: data = 8'b00000000;	//         
        11'h352: data = 8'b11111110;	// ******* 
        11'h353: data = 8'b11000000;	// **      
        11'h354: data = 8'b11000000;	// **      
        11'h355: data = 8'b01000000;	//  *      
        11'h356: data = 8'b00111100;	//   ****  
        11'h357: data = 8'b00000010;	//       * 
        11'h358: data = 8'b00000010;	//       * 
        11'h359: data = 8'b11111100;	// ******  
        11'h35a: data = 8'b00000000;	//         
        11'h35b: data = 8'b00000000;	//         
        11'h35c: data = 8'b00000000;	//         
        11'h35d: data = 8'b00000000;	//         
        11'h35e: data = 8'b00000000;	//         
        11'h35f: data = 8'b00000000;	//         

    // code x36 (6)
        11'h360: data = 8'b00000000;	//         
        11'h361: data = 8'b00000000;	//         
        11'h362: data = 8'b00111100;	//   ****  
        11'h363: data = 8'b00000010;	//       * 
        11'h364: data = 8'b11000000;	// **      
        11'h365: data = 8'b11000000;	// **      
        11'h366: data = 8'b11111100;	// ******  
        11'h367: data = 8'b11000010;	// **    * 
        11'h368: data = 8'b01000010;	//  *    * 
        11'h369: data = 8'b00111100;	//   ****  
        11'h36a: data = 8'b00000000;	//         
        11'h36b: data = 8'b00000000;	//         
        11'h36c: data = 8'b00000000;	//         
        11'h36d: data = 8'b00000000;	//         
        11'h36e: data = 8'b00000000;	//         
        11'h36f: data = 8'b00000000;	//         

    // code x37 (7)
        11'h370: data = 8'b00000000;	//         
        11'h371: data = 8'b00000000;	//         
        11'h372: data = 8'b11111100;	// ******  
        11'h373: data = 8'b00000010;	//       * 
        11'h374: data = 8'b00000010;	//       * 
        11'h375: data = 8'b00000010;	//       * 
        11'h376: data = 8'b00011110;	//    **** 
        11'h377: data = 8'b00000010;	//       * 
        11'h378: data = 8'b00000010;	//       * 
        11'h379: data = 8'b00000010;	//       * 
        11'h37a: data = 8'b00000000;	//         
        11'h37b: data = 8'b00000000;	//         
        11'h37c: data = 8'b00000000;	//         
        11'h37d: data = 8'b00000000;	//         
        11'h37e: data = 8'b00000000;	//         
        11'h37f: data = 8'b00000000;	//         

    // code x38 (8)
        11'h380: data = 8'b00000000;	//         
        11'h381: data = 8'b00000000;	//         
        11'h382: data = 8'b00111100;	//   ****  
        11'h383: data = 8'b11000010;	// **    * 
        11'h384: data = 8'b11000010;	// **    * 
        11'h385: data = 8'b00000000;	//         
        11'h386: data = 8'b00111100;	//   ****  
        11'h387: data = 8'b11000010;	// **    * 
        11'h388: data = 8'b11000010;	// **    * 
        11'h389: data = 8'b00111100;	//   ****  
        11'h38a: data = 8'b00000000;	//         
        11'h38b: data = 8'b00000000;	//         
        11'h38c: data = 8'b00000000;	//         
        11'h38d: data = 8'b00000000;	//         
        11'h38e: data = 8'b00000000;	//         
        11'h38f: data = 8'b00000000;	//         

    // code x39 (9)
        11'h390: data = 8'b00000000;	//         
        11'h391: data = 8'b00000000;	//         
        11'h392: data = 8'b00111100;	//   ****  
        11'h393: data = 8'b11000010;	// **    * 
        11'h394: data = 8'b11000010;	// **    * 
        11'h395: data = 8'b00000010;	//       * 
        11'h396: data = 8'b00111110;	//   ***** 
        11'h397: data = 8'b00000010;	//       * 
        11'h398: data = 8'b11000010;	// **    * 
        11'h399: data = 8'b00111100;	//   ****  
        11'h39a: data = 8'b00000000;	//         
        11'h39b: data = 8'b00000000;	//         
        11'h39c: data = 8'b00000000;	//         
        11'h39d: data = 8'b00000000;	//         
        11'h39e: data = 8'b00000000;	//         
        11'h39f: data = 8'b00000000;	//         

    // code xe01 (ก)
        11'he010: data = 8'b00000000;	//         
        11'he011: data = 8'b00000000;	//         
        11'he012: data = 8'b00000000;	//         
        11'he013: data = 8'b00111100;	//   ****  
        11'he014: data = 8'b11000010;	// **    * 
        11'he015: data = 8'b11000010;	// **    * 
        11'he016: data = 8'b11000010;	// **    * 
        11'he017: data = 8'b11000010;	// **    * 
        11'he018: data = 8'b11000010;	// **    * 
        11'he019: data = 8'b11000010;	// **    * 
        11'he01a: data = 8'b00000000;	//         
        11'he01b: data = 8'b00000000;	//         
        11'he01c: data = 8'b00000000;	//         
        11'he01d: data = 8'b00000000;	//         
        11'he01e: data = 8'b00000000;	//         
        11'he01f: data = 8'b00000000;	//         

    // code xe02 (ข)
        11'he020: data = 8'b00000000;	//         
        11'he021: data = 8'b00000000;	//         
        11'he022: data = 8'b00000000;	//         
        11'he023: data = 8'b11001000;	// **  *   
        11'he024: data = 8'b11001000;	// **  *   
        11'he025: data = 8'b11001000;	// **  *   
        11'he026: data = 8'b11001000;	// **  *   
        11'he027: data = 8'b11001000;	// **  *   
        11'he028: data = 8'b11001000;	// **  *   
        11'he029: data = 8'b00110000;	//   **    
        11'he02a: data = 8'b00000000;	//         
        11'he02b: data = 8'b00000000;	//         
        11'he02c: data = 8'b00000000;	//         
        11'he02d: data = 8'b00000000;	//         
        11'he02e: data = 8'b00000000;	//         
        11'he02f: data = 8'b00000000;	//         

    // code xe03 (ฃ)
        11'he030: data = 8'b00000000;	//         
        11'he031: data = 8'b00000000;	//         
        11'he032: data = 8'b00000000;	//         
        11'he033: data = 8'b10000100;	// *    *  
        11'he034: data = 8'b00100100;	//   *  *  
        11'he035: data = 8'b00100100;	//   *  *  
        11'he036: data = 8'b00100100;	//   *  *  
        11'he037: data = 8'b00100100;	//   *  *  
        11'he038: data = 8'b00100100;	//   *  *  
        11'he039: data = 8'b00011000;	//    **   
        11'he03a: data = 8'b00000000;	//         
        11'he03b: data = 8'b00000000;	//         
        11'he03c: data = 8'b00000000;	//         
        11'he03d: data = 8'b00000000;	//         
        11'he03e: data = 8'b00000000;	//         
        11'he03f: data = 8'b00000000;	//         

    // code xe04 (ค)
        11'he040: data = 8'b00000000;	//         
        11'he041: data = 8'b00000000;	//         
        11'he042: data = 8'b00000000;	//         
        11'he043: data = 8'b00111100;	//   ****  
        11'he044: data = 8'b11000010;	// **    * 
        11'he045: data = 8'b11000010;	// **    * 
        11'he046: data = 8'b11000010;	// **    * 
        11'he047: data = 8'b11110010;	// ****  * 
        11'he048: data = 8'b11000010;	// **    * 
        11'he049: data = 8'b11000010;	// **    * 
        11'he04a: data = 8'b00000000;	//         
        11'he04b: data = 8'b00000000;	//         
        11'he04c: data = 8'b00000000;	//         
        11'he04d: data = 8'b00000000;	//         
        11'he04e: data = 8'b00000000;	//         
        11'he04f: data = 8'b00000000;	//         

    // code xe05 (ฅ)
        11'he050: data = 8'b00000000;	//         
        11'he051: data = 8'b00000000;	//         
        11'he052: data = 8'b00000000;	//         
        11'he053: data = 8'b00100100;	//   *  *  
        11'he054: data = 8'b11000010;	// **    * 
        11'he055: data = 8'b11000010;	// **    * 
        11'he056: data = 8'b11000010;	// **    * 
        11'he057: data = 8'b11110010;	// ****  * 
        11'he058: data = 8'b11000010;	// **    * 
        11'he059: data = 8'b11000010;	// **    * 
        11'he05a: data = 8'b00000000;	//         
        11'he05b: data = 8'b00000000;	//         
        11'he05c: data = 8'b00000000;	//         
        11'he05d: data = 8'b00000000;	//         
        11'he05e: data = 8'b00000000;	//         
        11'he05f: data = 8'b00000000;	//         

    // code xe06 (ฆ)
        11'he060: data = 8'b00000000;	//         
        11'he061: data = 8'b00000000;	//         
        11'he062: data = 8'b00000000;	//         
        11'he063: data = 8'b10000010;	// *     * 
        11'he064: data = 8'b00100010;	//   *   * 
        11'he065: data = 8'b00100010;	//   *   * 
        11'he066: data = 8'b00100010;	//   *   * 
        11'he067: data = 8'b00100010;	//   *   * 
        11'he068: data = 8'b01110000;	//  ***    
        11'he069: data = 8'b00100100;	//   *  *  
        11'he06a: data = 8'b00000000;	//         
        11'he06b: data = 8'b00000000;	//         
        11'he06c: data = 8'b00000000;	//         
        11'he06d: data = 8'b00000000;	//         
        11'he06e: data = 8'b00000000;	//         
        11'he06f: data = 8'b00000000;	//         

    // code xe07 (ง)
        11'he070: data = 8'b00000000;	//         
        11'he071: data = 8'b00000000;	//         
        11'he072: data = 8'b00000000;	//         
        11'he073: data = 8'b00011000;	//    **   
        11'he074: data = 8'b00001000;	//     *   
        11'he075: data = 8'b00001000;	//     *   
        11'he076: data = 8'b11001000;	// **  *   
        11'he077: data = 8'b11001000;	// **  *   
        11'he078: data = 8'b11001000;	// **  *   
        11'he079: data = 8'b00110000;	//   **    
        11'he07a: data = 8'b00000000;	//         
        11'he07b: data = 8'b00000000;	//         
        11'he07c: data = 8'b00000000;	//         
        11'he07d: data = 8'b00000000;	//         
        11'he07e: data = 8'b00000000;	//         
        11'he07f: data = 8'b00000000;	//         

    // code xe08 (จ)
        11'he080: data = 8'b00000000;	//         
        11'he081: data = 8'b00000000;	//         
        11'he082: data = 8'b00000000;	//         
        11'he083: data = 8'b00111100;	//   ****  
        11'he084: data = 8'b00000010;	//       * 
        11'he085: data = 8'b11000010;	// **    * 
        11'he086: data = 8'b00000010;	//       * 
        11'he087: data = 8'b00001110;	//     *** 
        11'he088: data = 8'b00000010;	//       * 
        11'he089: data = 8'b00000010;	//       * 
        11'he08a: data = 8'b00000000;	//         
        11'he08b: data = 8'b00000000;	//         
        11'he08c: data = 8'b00000000;	//         
        11'he08d: data = 8'b00000000;	//         
        11'he08e: data = 8'b00000000;	//         
        11'he08f: data = 8'b00000000;	//         

    // code xe09 (ฉ)
        11'he090: data = 8'b00000000;	//         
        11'he091: data = 8'b00000000;	//         
        11'he092: data = 8'b00000000;	//         
        11'he093: data = 8'b00111100;	//   ****  
        11'he094: data = 8'b11000000;	// **      
        11'he095: data = 8'b11000010;	// **    * 
        11'he096: data = 8'b00000010;	//       * 
        11'he097: data = 8'b11000010;	// **    * 
        11'he098: data = 8'b11001111;	// **  ****
        11'he099: data = 8'b00100010;	//   *   * 
        11'he09a: data = 8'b00000000;	//         
        11'he09b: data = 8'b00000000;	//         
        11'he09c: data = 8'b00000000;	//         
        11'he09d: data = 8'b00000000;	//         
        11'he09e: data = 8'b00000000;	//         
        11'he09f: data = 8'b00000000;	//         

    // code xe0a (ช)
        11'he0a0: data = 8'b00000000;	//         
        11'he0a1: data = 8'b00000000;	//         
        11'he0a2: data = 8'b00000000;	//         
        11'he0a3: data = 8'b11001000;	// **  *   
        11'he0a4: data = 8'b11110000;	// ****    
        11'he0a5: data = 8'b11000000;	// **      
        11'he0a6: data = 8'b11001000;	// **  *   
        11'he0a7: data = 8'b11001000;	// **  *   
        11'he0a8: data = 8'b01001000;	//  *  *   
        11'he0a9: data = 8'b00110000;	//   **    
        11'he0aa: data = 8'b00000000;	//         
        11'he0ab: data = 8'b00000000;	//         
        11'he0ac: data = 8'b00000000;	//         
        11'he0ad: data = 8'b00000000;	//         
        11'he0ae: data = 8'b00000000;	//         
        11'he0af: data = 8'b00000000;	//         

    // code xe0b (ซ)
        11'he0b0: data = 8'b00000000;	//         
        11'he0b1: data = 8'b00000000;	//         
        11'he0b2: data = 8'b00000000;	//         
        11'he0b3: data = 8'b10000100;	// *    *  
        11'he0b4: data = 8'b00011000;	//    **   
        11'he0b5: data = 8'b00111000;	//   ***   
        11'he0b6: data = 8'b00100100;	//   *  *  
        11'he0b7: data = 8'b00100100;	//   *  *  
        11'he0b8: data = 8'b00100100;	//   *  *  
        11'he0b9: data = 8'b00011000;	//    **   
        11'he0ba: data = 8'b00000000;	//         
        11'he0bb: data = 8'b00000000;	//         
        11'he0bc: data = 8'b00000000;	//         
        11'he0bd: data = 8'b00000000;	//         
        11'he0be: data = 8'b00000000;	//         
        11'he0bf: data = 8'b00000000;	//         

    // code xe0c (ฌ)
        11'he0c0: data = 8'b00000000;	//         
        11'he0c1: data = 8'b00000000;	//         
        11'he0c2: data = 8'b00000000;	//         
        11'he0c3: data = 8'b00111100;	//   ****  
        11'he0c4: data = 8'b11000010;	// **    * 
        11'he0c5: data = 8'b11000010;	// **    * 
        11'he0c6: data = 8'b11000010;	// **    * 
        11'he0c7: data = 8'b11000010;	// **    * 
        11'he0c8: data = 8'b11000111;	// **   ***
        11'he0c9: data = 8'b11100010;	// ***   * 
        11'he0ca: data = 8'b00000000;	//         
        11'he0cb: data = 8'b00000000;	//         
        11'he0cc: data = 8'b00000000;	//         
        11'he0cd: data = 8'b00000000;	//         
        11'he0ce: data = 8'b00000000;	//         
        11'he0cf: data = 8'b00000000;	//         

    // code xe0d (ญ)
        11'he0d0: data = 8'b00000000;	//         
        11'he0d1: data = 8'b00000000;	//         
        11'he0d2: data = 8'b00000000;	//         
        11'he0d3: data = 8'b00111100;	//   ****  
        11'he0d4: data = 8'b11000010;	// **    * 
        11'he0d5: data = 8'b11000010;	// **    * 
        11'he0d6: data = 8'b11000010;	// **    * 
        11'he0d7: data = 8'b11000010;	// **    * 
        11'he0d8: data = 8'b11000001;	// **     *
        11'he0d9: data = 8'b11100000;	// ***     
        11'he0da: data = 8'b00000001;	//        *
        11'he0db: data = 8'b00000000;	//         
        11'he0dc: data = 8'b00000000;	//         
        11'he0dd: data = 8'b00000000;	//         
        11'he0de: data = 8'b00000000;	//         
        11'he0df: data = 8'b00000000;	//         

    // code xe0e (ฎ)
        11'he0e0: data = 8'b00000000;	//         
        11'he0e1: data = 8'b00000000;	//         
        11'he0e2: data = 8'b00000000;	//         
        11'he0e3: data = 8'b00111100;	//   ****  
        11'he0e4: data = 8'b11000010;	// **    * 
        11'he0e5: data = 8'b11000010;	// **    * 
        11'he0e6: data = 8'b11000010;	// **    * 
        11'he0e7: data = 8'b11000010;	// **    * 
        11'he0e8: data = 8'b11000010;	// **    * 
        11'he0e9: data = 8'b11000010;	// **    * 
        11'he0ea: data = 8'b00000010;	//       * 
        11'he0eb: data = 8'b00100100;	//   *  *  
        11'he0ec: data = 8'b00000000;	//         
        11'he0ed: data = 8'b00000000;	//         
        11'he0ee: data = 8'b00000000;	//         
        11'he0ef: data = 8'b00000000;	//         

    // code xe0f (ฏ)
        11'he0f0: data = 8'b00000000;	//         
        11'he0f1: data = 8'b00000000;	//         
        11'he0f2: data = 8'b00000000;	//         
        11'he0f3: data = 8'b00111100;	//   ****  
        11'he0f4: data = 8'b11000010;	// **    * 
        11'he0f5: data = 8'b11000010;	// **    * 
        11'he0f6: data = 8'b11000010;	// **    * 
        11'he0f7: data = 8'b11000010;	// **    * 
        11'he0f8: data = 8'b11000010;	// **    * 
        11'he0f9: data = 8'b11000010;	// **    * 
        11'he0fa: data = 8'b00000110;	//      ** 
        11'he0fb: data = 8'b00000010;	//       * 
        11'he0fc: data = 8'b00000000;	//         
        11'he0fd: data = 8'b00000000;	//         
        11'he0fe: data = 8'b00000000;	//         
        11'he0ff: data = 8'b00000000;	//         

    // code xe10 (ฐ)
        11'he100: data = 8'b00000000;	//         
        11'he101: data = 8'b00000000;	//         
        11'he102: data = 8'b00000000;	//         
        11'he103: data = 8'b00111110;	//   ***** 
        11'he104: data = 8'b00000010;	//       * 
        11'he105: data = 8'b00000010;	//       * 
        11'he106: data = 8'b00000010;	//       * 
        11'he107: data = 8'b00001110;	//     *** 
        11'he108: data = 8'b00000010;	//       * 
        11'he109: data = 8'b00000010;	//       * 
        11'he10a: data = 8'b00000000;	//         
        11'he10b: data = 8'b00000000;	//         
        11'he10c: data = 8'b00000000;	//         
        11'he10d: data = 8'b00000000;	//         
        11'he10e: data = 8'b00000000;	//         
        11'he10f: data = 8'b00000000;	//         

    // code xe11 (ฑ)
        11'he110: data = 8'b00000000;	//         
        11'he111: data = 8'b00000000;	//         
        11'he112: data = 8'b00000000;	//         
        11'he113: data = 8'b10000010;	// *     * 
        11'he114: data = 8'b00100001;	//   *    *
        11'he115: data = 8'b00100001;	//   *    *
        11'he116: data = 8'b00110001;	//   **   *
        11'he117: data = 8'b00100001;	//   *    *
        11'he118: data = 8'b00100001;	//   *    *
        11'he119: data = 8'b00100001;	//   *    *
        11'he11a: data = 8'b00000000;	//         
        11'he11b: data = 8'b00000000;	//         
        11'he11c: data = 8'b00000000;	//         
        11'he11d: data = 8'b00000000;	//         
        11'he11e: data = 8'b00000000;	//         
        11'he11f: data = 8'b00000000;	//         

    // code xe12 (ฒ)
        11'he120: data = 8'b00000000;	//         
        11'he121: data = 8'b00000000;	//         
        11'he122: data = 8'b00000000;	//         
        11'he123: data = 8'b00100100;	//   *  *  
        11'he124: data = 8'b11000010;	// **    * 
        11'he125: data = 8'b11000010;	// **    * 
        11'he126: data = 8'b11000010;	// **    * 
        11'he127: data = 8'b11000010;	// **    * 
        11'he128: data = 8'b11000111;	// **   ***
        11'he129: data = 8'b00100010;	//   *   * 
        11'he12a: data = 8'b00000000;	//         
        11'he12b: data = 8'b00000000;	//         
        11'he12c: data = 8'b00000000;	//         
        11'he12d: data = 8'b00000000;	//         
        11'he12e: data = 8'b00000000;	//         
        11'he12f: data = 8'b00000000;	//         

    // code xe13 (ณ)
        11'he130: data = 8'b00000000;	//         
        11'he131: data = 8'b00000000;	//         
        11'he132: data = 8'b00000000;	//         
        11'he133: data = 8'b00111100;	//   ****  
        11'he134: data = 8'b11000010;	// **    * 
        11'he135: data = 8'b11000010;	// **    * 
        11'he136: data = 8'b11000010;	// **    * 
        11'he137: data = 8'b11000010;	// **    * 
        11'he138: data = 8'b11000010;	// **    * 
        11'he139: data = 8'b11100001;	// ***    *
        11'he13a: data = 8'b00000000;	//         
        11'he13b: data = 8'b00000000;	//         
        11'he13c: data = 8'b00000000;	//         
        11'he13d: data = 8'b00000000;	//         
        11'he13e: data = 8'b00000000;	//         
        11'he13f: data = 8'b00000000;	//         

    // code xe14 (ด)
        11'he140: data = 8'b00000000;	//         
        11'he141: data = 8'b00000000;	//         
        11'he142: data = 8'b00000000;	//         
        11'he143: data = 8'b00111100;	//   ****  
        11'he144: data = 8'b11000010;	// **    * 
        11'he145: data = 8'b11000010;	// **    * 
        11'he146: data = 8'b11000010;	// **    * 
        11'he147: data = 8'b11000010;	// **    * 
        11'he148: data = 8'b11000010;	// **    * 
        11'he149: data = 8'b00110010;	//   **  * 
        11'he14a: data = 8'b00000000;	//         
        11'he14b: data = 8'b00000000;	//         
        11'he14c: data = 8'b00000000;	//         
        11'he14d: data = 8'b00000000;	//         
        11'he14e: data = 8'b00000000;	//         
        11'he14f: data = 8'b00000000;	//         

    // code xe15 (ต)
        11'he150: data = 8'b00000000;	//         
        11'he151: data = 8'b00000000;	//         
        11'he152: data = 8'b00000000;	//         
        11'he153: data = 8'b00100100;	//   *  *  
        11'he154: data = 8'b11000010;	// **    * 
        11'he155: data = 8'b11000010;	// **    * 
        11'he156: data = 8'b11000010;	// **    * 
        11'he157: data = 8'b11000010;	// **    * 
        11'he158: data = 8'b11000010;	// **    * 
        11'he159: data = 8'b00110010;	//   **  * 
        11'he15a: data = 8'b00000000;	//         
        11'he15b: data = 8'b00000000;	//         
        11'he15c: data = 8'b00000000;	//         
        11'he15d: data = 8'b00000000;	//         
        11'he15e: data = 8'b00000000;	//         
        11'he15f: data = 8'b00000000;	//         

    // code xe16 (ถ)
        11'he160: data = 8'b00000000;	//         
        11'he161: data = 8'b00000000;	//         
        11'he162: data = 8'b00000000;	//         
        11'he163: data = 8'b00111100;	//   ****  
        11'he164: data = 8'b11000010;	// **    * 
        11'he165: data = 8'b11000010;	// **    * 
        11'he166: data = 8'b11000010;	// **    * 
        11'he167: data = 8'b11000010;	// **    * 
        11'he168: data = 8'b11000010;	// **    * 
        11'he169: data = 8'b11100010;	// ***   * 
        11'he16a: data = 8'b00000000;	//         
        11'he16b: data = 8'b00000000;	//         
        11'he16c: data = 8'b00000000;	//         
        11'he16d: data = 8'b00000000;	//         
        11'he16e: data = 8'b00000000;	//         
        11'he16f: data = 8'b00000000;	//         

    // code xe17 (ท)
        11'he170: data = 8'b00000000;	//         
        11'he171: data = 8'b00000000;	//         
        11'he172: data = 8'b00000000;	//         
        11'he173: data = 8'b11000100;	// **   *  
        11'he174: data = 8'b11000010;	// **    * 
        11'he175: data = 8'b11100010;	// ***   * 
        11'he176: data = 8'b11000010;	// **    * 
        11'he177: data = 8'b11000010;	// **    * 
        11'he178: data = 8'b11000010;	// **    * 
        11'he179: data = 8'b11000010;	// **    * 
        11'he17a: data = 8'b00000000;	//         
        11'he17b: data = 8'b00000000;	//         
        11'he17c: data = 8'b00000000;	//         
        11'he17d: data = 8'b00000000;	//         
        11'he17e: data = 8'b00000000;	//         
        11'he17f: data = 8'b00000000;	//         

    // code xe18 (ธ)
        11'he180: data = 8'b00000000;	//         
        11'he181: data = 8'b00000000;	//         
        11'he182: data = 8'b00000000;	//         
        11'he183: data = 8'b00111110;	//   ***** 
        11'he184: data = 8'b11000000;	// **      
        11'he185: data = 8'b00000000;	//         
        11'he186: data = 8'b00111100;	//   ****  
        11'he187: data = 8'b00000010;	//       * 
        11'he188: data = 8'b11000010;	// **    * 
        11'he189: data = 8'b11111100;	// ******  
        11'he18a: data = 8'b00000000;	//         
        11'he18b: data = 8'b00000000;	//         
        11'he18c: data = 8'b00000000;	//         
        11'he18d: data = 8'b00000000;	//         
        11'he18e: data = 8'b00000000;	//         
        11'he18f: data = 8'b00000000;	//         

    // code xe19 (น)
        11'he190: data = 8'b00000000;	//         
        11'he191: data = 8'b00000000;	//         
        11'he192: data = 8'b00000000;	//         
        11'he193: data = 8'b11000010;	// **    * 
        11'he194: data = 8'b11000010;	// **    * 
        11'he195: data = 8'b11000010;	// **    * 
        11'he196: data = 8'b11000010;	// **    * 
        11'he197: data = 8'b11000010;	// **    * 
        11'he198: data = 8'b01000011;	//  *    **
        11'he199: data = 8'b00100010;	//   *   * 
        11'he19a: data = 8'b00000000;	//         
        11'he19b: data = 8'b00000000;	//         
        11'he19c: data = 8'b00000000;	//         
        11'he19d: data = 8'b00000000;	//         
        11'he19e: data = 8'b00000000;	//         
        11'he19f: data = 8'b00000000;	//         

    // code xe1a (บ)
        11'he1a0: data = 8'b00000000;	//         
        11'he1a1: data = 8'b00000000;	//         
        11'he1a2: data = 8'b00000000;	//         
        11'he1a3: data = 8'b11000010;	// **    * 
        11'he1a4: data = 8'b11000010;	// **    * 
        11'he1a5: data = 8'b11000010;	// **    * 
        11'he1a6: data = 8'b11000010;	// **    * 
        11'he1a7: data = 8'b11000010;	// **    * 
        11'he1a8: data = 8'b11000010;	// **    * 
        11'he1a9: data = 8'b00111100;	//   ****  
        11'he1aa: data = 8'b00000000;	//         
        11'he1ab: data = 8'b00000000;	//         
        11'he1ac: data = 8'b00000000;	//         
        11'he1ad: data = 8'b00000000;	//         
        11'he1ae: data = 8'b00000000;	//         
        11'he1af: data = 8'b00000000;	//         

    // code xe1b (ป)
        11'he1b0: data = 8'b00000000;	//         
        11'he1b1: data = 8'b00000010;	//       * 
        11'he1b2: data = 8'b00000010;	//       * 
        11'he1b3: data = 8'b00000010;	//       * 
        11'he1b4: data = 8'b11000010;	// **    * 
        11'he1b5: data = 8'b11000010;	// **    * 
        11'he1b6: data = 8'b11000010;	// **    * 
        11'he1b7: data = 8'b11000010;	// **    * 
        11'he1b8: data = 8'b11000010;	// **    * 
        11'he1b9: data = 8'b00111100;	//   ****  
        11'he1ba: data = 8'b00000000;	//         
        11'he1bb: data = 8'b00000000;	//         
        11'he1bc: data = 8'b00000000;	//         
        11'he1bd: data = 8'b00000000;	//         
        11'he1be: data = 8'b00000000;	//         
        11'he1bf: data = 8'b00000000;	//         

    // code xe1c (ผ)
        11'he1c0: data = 8'b00000000;	//         
        11'he1c1: data = 8'b00000000;	//         
        11'he1c2: data = 8'b00000000;	//         
        11'he1c3: data = 8'b00100010;	//   *   * 
        11'he1c4: data = 8'b11000010;	// **    * 
        11'he1c5: data = 8'b11000010;	// **    * 
        11'he1c6: data = 8'b11000010;	// **    * 
        11'he1c7: data = 8'b11000010;	// **    * 
        11'he1c8: data = 8'b11000010;	// **    * 
        11'he1c9: data = 8'b00100100;	//   *  *  
        11'he1ca: data = 8'b00000000;	//         
        11'he1cb: data = 8'b00000000;	//         
        11'he1cc: data = 8'b00000000;	//         
        11'he1cd: data = 8'b00000000;	//         
        11'he1ce: data = 8'b00000000;	//         
        11'he1cf: data = 8'b00000000;	//         

    // code xe1d (ฝ)
        11'he1d0: data = 8'b00000000;	//         
        11'he1d1: data = 8'b00000010;	//       * 
        11'he1d2: data = 8'b00000010;	//       * 
        11'he1d3: data = 8'b00100010;	//   *   * 
        11'he1d4: data = 8'b11000010;	// **    * 
        11'he1d5: data = 8'b11000010;	// **    * 
        11'he1d6: data = 8'b11000010;	// **    * 
        11'he1d7: data = 8'b11000010;	// **    * 
        11'he1d8: data = 8'b11000010;	// **    * 
        11'he1d9: data = 8'b00100100;	//   *  *  
        11'he1da: data = 8'b00000000;	//         
        11'he1db: data = 8'b00000000;	//         
        11'he1dc: data = 8'b00000000;	//         
        11'he1dd: data = 8'b00000000;	//         
        11'he1de: data = 8'b00000000;	//         
        11'he1df: data = 8'b00000000;	//         

    // code xe1e (พ)
        11'he1e0: data = 8'b00000000;	//         
        11'he1e1: data = 8'b00000000;	//         
        11'he1e2: data = 8'b00000000;	//         
        11'he1e3: data = 8'b11000010;	// **    * 
        11'he1e4: data = 8'b11000010;	// **    * 
        11'he1e5: data = 8'b11000010;	// **    * 
        11'he1e6: data = 8'b11000010;	// **    * 
        11'he1e7: data = 8'b11000010;	// **    * 
        11'he1e8: data = 8'b11000010;	// **    * 
        11'he1e9: data = 8'b00100100;	//   *  *  
        11'he1ea: data = 8'b00000000;	//         
        11'he1eb: data = 8'b00000000;	//         
        11'he1ec: data = 8'b00000000;	//         
        11'he1ed: data = 8'b00000000;	//         
        11'he1ee: data = 8'b00000000;	//         
        11'he1ef: data = 8'b00000000;	//         

    // code xe1f (ฟ)
        11'he1f0: data = 8'b00000000;	//         
        11'he1f1: data = 8'b00000010;	//       * 
        11'he1f2: data = 8'b00000010;	//       * 
        11'he1f3: data = 8'b00000010;	//       * 
        11'he1f4: data = 8'b11000010;	// **    * 
        11'he1f5: data = 8'b11000010;	// **    * 
        11'he1f6: data = 8'b11000010;	// **    * 
        11'he1f7: data = 8'b11000010;	// **    * 
        11'he1f8: data = 8'b11000010;	// **    * 
        11'he1f9: data = 8'b00100100;	//   *  *  
        11'he1fa: data = 8'b00000000;	//         
        11'he1fb: data = 8'b00000000;	//         
        11'he1fc: data = 8'b00000000;	//         
        11'he1fd: data = 8'b00000000;	//         
        11'he1fe: data = 8'b00000000;	//         
        11'he1ff: data = 8'b00000000;	//         

    // code xe20 (ภ)
        11'he200: data = 8'b00000000;	//         
        11'he201: data = 8'b00000000;	//         
        11'he202: data = 8'b00000000;	//         
        11'he203: data = 8'b00011110;	//    **** 
        11'he204: data = 8'b00100001;	//   *    *
        11'he205: data = 8'b00100001;	//   *    *
        11'he206: data = 8'b00100001;	//   *    *
        11'he207: data = 8'b00100001;	//   *    *
        11'he208: data = 8'b00100001;	//   *    *
        11'he209: data = 8'b11100001;	// ***    *
        11'he20a: data = 8'b00000000;	//         
        11'he20b: data = 8'b00000000;	//         
        11'he20c: data = 8'b00000000;	//         
        11'he20d: data = 8'b00000000;	//         
        11'he20e: data = 8'b00000000;	//         
        11'he20f: data = 8'b00000000;	//         

    // code xe21 (ม)
        11'he210: data = 8'b00000000;	//         
        11'he211: data = 8'b00000000;	//         
        11'he212: data = 8'b00000000;	//         
        11'he213: data = 8'b11100001;	// ***    *
        11'he214: data = 8'b00100001;	//   *    *
        11'he215: data = 8'b00100001;	//   *    *
        11'he216: data = 8'b00100001;	//   *    *
        11'he217: data = 8'b00100001;	//   *    *
        11'he218: data = 8'b11111001;	// *****  *
        11'he219: data = 8'b00100010;	//   *   * 
        11'he21a: data = 8'b00000000;	//         
        11'he21b: data = 8'b00000000;	//         
        11'he21c: data = 8'b00000000;	//         
        11'he21d: data = 8'b00000000;	//         
        11'he21e: data = 8'b00000000;	//         
        11'he21f: data = 8'b00000000;	//         

    // code xe22 (ย)
        11'he220: data = 8'b00000000;	//         
        11'he221: data = 8'b00000000;	//         
        11'he222: data = 8'b00000000;	//         
        11'he223: data = 8'b00100010;	//   *   * 
        11'he224: data = 8'b11000010;	// **    * 
        11'he225: data = 8'b00000010;	//       * 
        11'he226: data = 8'b00110010;	//   **  * 
        11'he227: data = 8'b11000010;	// **    * 
        11'he228: data = 8'b11000010;	// **    * 
        11'he229: data = 8'b00111100;	//   ****  
        11'he22a: data = 8'b00000000;	//         
        11'he22b: data = 8'b00000000;	//         
        11'he22c: data = 8'b00000000;	//         
        11'he22d: data = 8'b00000000;	//         
        11'he22e: data = 8'b00000000;	//         
        11'he22f: data = 8'b00000000;	//         

    // code xe23 (ร)
        11'he230: data = 8'b00000000;	//         
        11'he231: data = 8'b00000000;	//         
        11'he232: data = 8'b00000000;	//         
        11'he233: data = 8'b00111100;	//   ****  
        11'he234: data = 8'b11000000;	// **      
        11'he235: data = 8'b00000000;	//         
        11'he236: data = 8'b00111000;	//   ***   
        11'he237: data = 8'b00000100;	//      *  
        11'he238: data = 8'b00000100;	//      *  
        11'he239: data = 8'b00011000;	//    **   
        11'he23a: data = 8'b00000000;	//         
        11'he23b: data = 8'b00000000;	//         
        11'he23c: data = 8'b00000000;	//         
        11'he23d: data = 8'b00000000;	//         
        11'he23e: data = 8'b00000000;	//         
        11'he23f: data = 8'b00000000;	//         

    // code xe24 (ฤ)
        11'he240: data = 8'b00000000;	//         
        11'he241: data = 8'b00000000;	//         
        11'he242: data = 8'b00000000;	//         
        11'he243: data = 8'b00111100;	//   ****  
        11'he244: data = 8'b11000010;	// **    * 
        11'he245: data = 8'b11000010;	// **    * 
        11'he246: data = 8'b11000010;	// **    * 
        11'he247: data = 8'b11000010;	// **    * 
        11'he248: data = 8'b11000010;	// **    * 
        11'he249: data = 8'b11100010;	// ***   * 
        11'he24a: data = 8'b00000010;	//       * 
        11'he24b: data = 8'b00000010;	//       * 
        11'he24c: data = 8'b00000000;	//         
        11'he24d: data = 8'b00000000;	//         
        11'he24e: data = 8'b00000000;	//         
        11'he24f: data = 8'b00000000;	//         

    // code xe25 (ล)
        11'he250: data = 8'b00000000;	//         
        11'he251: data = 8'b00000000;	//         
        11'he252: data = 8'b00000000;	//         
        11'he253: data = 8'b11111100;	// ******  
        11'he254: data = 8'b00000010;	//       * 
        11'he255: data = 8'b00000010;	//       * 
        11'he256: data = 8'b00111110;	//   ***** 
        11'he257: data = 8'b11000010;	// **    * 
        11'he258: data = 8'b01000010;	//  *    * 
        11'he259: data = 8'b00100010;	//   *   * 
        11'he25a: data = 8'b00000000;	//         
        11'he25b: data = 8'b00000000;	//         
        11'he25c: data = 8'b00000000;	//         
        11'he25d: data = 8'b00000000;	//         
        11'he25e: data = 8'b00000000;	//         
        11'he25f: data = 8'b00000000;	//         

    // code xe26 (ฦ)
        11'he260: data = 8'b00000000;	//         
        11'he261: data = 8'b00000000;	//         
        11'he262: data = 8'b00000000;	//         
        11'he263: data = 8'b00011110;	//    **** 
        11'he264: data = 8'b00100001;	//   *    *
        11'he265: data = 8'b00100001;	//   *    *
        11'he266: data = 8'b00100001;	//   *    *
        11'he267: data = 8'b00100001;	//   *    *
        11'he268: data = 8'b00100001;	//   *    *
        11'he269: data = 8'b11100001;	// ***    *
        11'he26a: data = 8'b00000001;	//        *
        11'he26b: data = 8'b00000001;	//        *
        11'he26c: data = 8'b00000000;	//         
        11'he26d: data = 8'b00000000;	//         
        11'he26e: data = 8'b00000000;	//         
        11'he26f: data = 8'b00000000;	//         

    // code xe27 (ว)
        11'he270: data = 8'b00000000;	//         
        11'he271: data = 8'b00000000;	//         
        11'he272: data = 8'b00000000;	//         
        11'he273: data = 8'b11111000;	// *****   
        11'he274: data = 8'b00000100;	//      *  
        11'he275: data = 8'b00000100;	//      *  
        11'he276: data = 8'b00000100;	//      *  
        11'he277: data = 8'b00000100;	//      *  
        11'he278: data = 8'b00000100;	//      *  
        11'he279: data = 8'b00011000;	//    **   
        11'he27a: data = 8'b00000000;	//         
        11'he27b: data = 8'b00000000;	//         
        11'he27c: data = 8'b00000000;	//         
        11'he27d: data = 8'b00000000;	//         
        11'he27e: data = 8'b00000000;	//         
        11'he27f: data = 8'b00000000;	//         

    // code xe28 (ศ)
        11'he280: data = 8'b00000000;	//         
        11'he281: data = 8'b00000000;	//         
        11'he282: data = 8'b00000010;	//       * 
        11'he283: data = 8'b00111110;	//   ***** 
        11'he284: data = 8'b11000010;	// **    * 
        11'he285: data = 8'b11000010;	// **    * 
        11'he286: data = 8'b11000010;	// **    * 
        11'he287: data = 8'b11110010;	// ****  * 
        11'he288: data = 8'b11000010;	// **    * 
        11'he289: data = 8'b11000010;	// **    * 
        11'he28a: data = 8'b00000000;	//         
        11'he28b: data = 8'b00000000;	//         
        11'he28c: data = 8'b00000000;	//         
        11'he28d: data = 8'b00000000;	//         
        11'he28e: data = 8'b00000000;	//         
        11'he28f: data = 8'b00000000;	//         

    // code xe29 (ษ)
        11'he290: data = 8'b00000000;	//         
        11'he291: data = 8'b00000000;	//         
        11'he292: data = 8'b00000000;	//         
        11'he293: data = 8'b11000010;	// **    * 
        11'he294: data = 8'b11000010;	// **    * 
        11'he295: data = 8'b11000010;	// **    * 
        11'he296: data = 8'b11001110;	// **  *** 
        11'he297: data = 8'b11000010;	// **    * 
        11'he298: data = 8'b11000010;	// **    * 
        11'he299: data = 8'b00111100;	//   ****  
        11'he29a: data = 8'b00000000;	//         
        11'he29b: data = 8'b00000000;	//         
        11'he29c: data = 8'b00000000;	//         
        11'he29d: data = 8'b00000000;	//         
        11'he29e: data = 8'b00000000;	//         
        11'he29f: data = 8'b00000000;	//         

    // code xe2a (ส)
        11'he2a0: data = 8'b00000000;	//         
        11'he2a1: data = 8'b00000000;	//         
        11'he2a2: data = 8'b00000010;	//       * 
        11'he2a3: data = 8'b11111110;	// ******* 
        11'he2a4: data = 8'b00000010;	//       * 
        11'he2a5: data = 8'b00000010;	//       * 
        11'he2a6: data = 8'b00111110;	//   ***** 
        11'he2a7: data = 8'b11000010;	// **    * 
        11'he2a8: data = 8'b01000010;	//  *    * 
        11'he2a9: data = 8'b00100010;	//   *   * 
        11'he2aa: data = 8'b00000000;	//         
        11'he2ab: data = 8'b00000000;	//         
        11'he2ac: data = 8'b00000000;	//         
        11'he2ad: data = 8'b00000000;	//         
        11'he2ae: data = 8'b00000000;	//         
        11'he2af: data = 8'b00000000;	//         

    // code xe2b (ห)
        11'he2b0: data = 8'b00000000;	//         
        11'he2b1: data = 8'b00000000;	//         
        11'he2b2: data = 8'b00000000;	//         
        11'he2b3: data = 8'b00000000;	//         
        11'he2b4: data = 8'b11000010;	// **    * 
        11'he2b5: data = 8'b11000010;	// **    * 
        11'he2b6: data = 8'b11000100;	// **   *  
        11'he2b7: data = 8'b11000010;	// **    * 
        11'he2b8: data = 8'b11100010;	// ***   * 
        11'he2b9: data = 8'b11000010;	// **    * 
        11'he2ba: data = 8'b00000000;	//         
        11'he2bb: data = 8'b00000000;	//         
        11'he2bc: data = 8'b00000000;	//         
        11'he2bd: data = 8'b00000000;	//         
        11'he2be: data = 8'b00000000;	//         
        11'he2bf: data = 8'b00000000;	//         

    // code xe2c (ฬ)
        11'he2c0: data = 8'b00000000;	//         
        11'he2c1: data = 8'b00000000;	//         
        11'he2c2: data = 8'b00000000;	//         
        11'he2c3: data = 8'b11000010;	// **    * 
        11'he2c4: data = 8'b11000100;	// **   *  
        11'he2c5: data = 8'b11000100;	// **   *  
        11'he2c6: data = 8'b11000010;	// **    * 
        11'he2c7: data = 8'b11000010;	// **    * 
        11'he2c8: data = 8'b01000010;	//  *    * 
        11'he2c9: data = 8'b00100100;	//   *  *  
        11'he2ca: data = 8'b00000000;	//         
        11'he2cb: data = 8'b00000000;	//         
        11'he2cc: data = 8'b00000000;	//         
        11'he2cd: data = 8'b00000000;	//         
        11'he2ce: data = 8'b00000000;	//         
        11'he2cf: data = 8'b00000000;	//         

    // code xe2d (อ)
        11'he2d0: data = 8'b00000000;	//         
        11'he2d1: data = 8'b00000000;	//         
        11'he2d2: data = 8'b00000000;	//         
        11'he2d3: data = 8'b11111100;	// ******  
        11'he2d4: data = 8'b00000010;	//       * 
        11'he2d5: data = 8'b00000010;	//       * 
        11'he2d6: data = 8'b11100010;	// ***   * 
        11'he2d7: data = 8'b11000010;	// **    * 
        11'he2d8: data = 8'b11000010;	// **    * 
        11'he2d9: data = 8'b00111100;	//   ****  
        11'he2da: data = 8'b00000000;	//         
        11'he2db: data = 8'b00000000;	//         
        11'he2dc: data = 8'b00000000;	//         
        11'he2dd: data = 8'b00000000;	//         
        11'he2de: data = 8'b00000000;	//         
        11'he2df: data = 8'b00000000;	//         

    // code xe2e (ฮ)
        11'he2e0: data = 8'b00000000;	//         
        11'he2e1: data = 8'b00000000;	//         
        11'he2e2: data = 8'b00000010;	//       * 
        11'he2e3: data = 8'b11111110;	// ******* 
        11'he2e4: data = 8'b00000010;	//       * 
        11'he2e5: data = 8'b00000010;	//       * 
        11'he2e6: data = 8'b11100010;	// ***   * 
        11'he2e7: data = 8'b11000010;	// **    * 
        11'he2e8: data = 8'b11000010;	// **    * 
        11'he2e9: data = 8'b00111100;	//   ****  
        11'he2ea: data = 8'b00000000;	//         
        11'he2eb: data = 8'b00000000;	//         
        11'he2ec: data = 8'b00000000;	//         
        11'he2ed: data = 8'b00000000;	//         
        11'he2ee: data = 8'b00000000;	//         
        11'he2ef: data = 8'b00000000;	//         

    // code xe2f (ฯ)
        11'he2f0: data = 8'b00000000;	//         
        11'he2f1: data = 8'b00000000;	//         
        11'he2f2: data = 8'b00000000;	//         
        11'he2f3: data = 8'b00100010;	//   *   * 
        11'he2f4: data = 8'b11000110;	// **   ** 
        11'he2f5: data = 8'b00110010;	//   **  * 
        11'he2f6: data = 8'b00110010;	//   **  * 
        11'he2f7: data = 8'b00000010;	//       * 
        11'he2f8: data = 8'b00000010;	//       * 
        11'he2f9: data = 8'b00011100;	//    ***  
        11'he2fa: data = 8'b00000000;	//         
        11'he2fb: data = 8'b00000000;	//         
        11'he2fc: data = 8'b00000000;	//         
        11'he2fd: data = 8'b00000000;	//         
        11'he2fe: data = 8'b00000000;	//         
        11'he2ff: data = 8'b00000000;	//         

    // code xe30 (ะ)
        11'he300: data = 8'b00000000;	//         
        11'he301: data = 8'b00000000;	//         
        11'he302: data = 8'b00000000;	//         
        11'he303: data = 8'b00000000;	//         
        11'he304: data = 8'b00000000;	//         
        11'he305: data = 8'b11000000;	// **      
        11'he306: data = 8'b11110000;	// ****    
        11'he307: data = 8'b00000000;	//         
        11'he308: data = 8'b11000000;	// **      
        11'he309: data = 8'b11110000;	// ****    
        11'he30a: data = 8'b00000000;	//         
        11'he30b: data = 8'b00000000;	//         
        11'he30c: data = 8'b00000000;	//         
        11'he30d: data = 8'b00000000;	//         
        11'he30e: data = 8'b00000000;	//         
        11'he30f: data = 8'b00000000;	//         

    // code xe31 (ั)
        11'he310: data = 8'b00000000;	//         
        11'he311: data = 8'b00000000;	//         
        11'he312: data = 8'b00000000;	//         
        11'he313: data = 8'b00000100;	//      *  
        11'he314: data = 8'b00000111;	//      ***
        11'he315: data = 8'b00000000;	//         
        11'he316: data = 8'b00000000;	//         
        11'he317: data = 8'b00000000;	//         
        11'he318: data = 8'b00000000;	//         
        11'he319: data = 8'b00000000;	//         
        11'he31a: data = 8'b00000000;	//         
        11'he31b: data = 8'b00000000;	//         
        11'he31c: data = 8'b00000000;	//         
        11'he31d: data = 8'b00000000;	//         
        11'he31e: data = 8'b00000000;	//         
        11'he31f: data = 8'b00000000;	//         

    // code xe32 (า)
        11'he320: data = 8'b00000000;	//         
        11'he321: data = 8'b00000000;	//         
        11'he322: data = 8'b00000000;	//         
        11'he323: data = 8'b11111000;	// *****   
        11'he324: data = 8'b00000100;	//      *  
        11'he325: data = 8'b00000100;	//      *  
        11'he326: data = 8'b00000100;	//      *  
        11'he327: data = 8'b00000100;	//      *  
        11'he328: data = 8'b00000100;	//      *  
        11'he329: data = 8'b00000100;	//      *  
        11'he32a: data = 8'b00000000;	//         
        11'he32b: data = 8'b00000000;	//         
        11'he32c: data = 8'b00000000;	//         
        11'he32d: data = 8'b00000000;	//         
        11'he32e: data = 8'b00000000;	//         
        11'he32f: data = 8'b00000000;	//         

    // code xe33 (ำ)
        11'he330: data = 8'b00000000;	//         
        11'he331: data = 8'b00000000;	//         
        11'he332: data = 8'b00000000;	//         
        11'he333: data = 8'b11111000;	// *****   
        11'he334: data = 8'b00000100;	//      *  
        11'he335: data = 8'b00000100;	//      *  
        11'he336: data = 8'b00000100;	//      *  
        11'he337: data = 8'b00000100;	//      *  
        11'he338: data = 8'b00000100;	//      *  
        11'he339: data = 8'b00000100;	//      *  
        11'he33a: data = 8'b00000000;	//         
        11'he33b: data = 8'b00000000;	//         
        11'he33c: data = 8'b00000000;	//         
        11'he33d: data = 8'b00000000;	//         
        11'he33e: data = 8'b00000000;	//         
        11'he33f: data = 8'b00000000;	//         

    // code xe34 (ิ)
        11'he340: data = 8'b00000000;	//         
        11'he341: data = 8'b00000000;	//         
        11'he342: data = 8'b00000000;	//         
        11'he343: data = 8'b00000000;	//         
        11'he344: data = 8'b00001111;	//     ****
        11'he345: data = 8'b00000000;	//         
        11'he346: data = 8'b00000000;	//         
        11'he347: data = 8'b00000000;	//         
        11'he348: data = 8'b00000000;	//         
        11'he349: data = 8'b00000000;	//         
        11'he34a: data = 8'b00000000;	//         
        11'he34b: data = 8'b00000000;	//         
        11'he34c: data = 8'b00000000;	//         
        11'he34d: data = 8'b00000000;	//         
        11'he34e: data = 8'b00000000;	//         
        11'he34f: data = 8'b00000000;	//         

    // code xe35 (ี)
        11'he350: data = 8'b00000000;	//         
        11'he351: data = 8'b00000000;	//         
        11'he352: data = 8'b00000000;	//         
        11'he353: data = 8'b00000001;	//        *
        11'he354: data = 8'b00001111;	//     ****
        11'he355: data = 8'b00000000;	//         
        11'he356: data = 8'b00000000;	//         
        11'he357: data = 8'b00000000;	//         
        11'he358: data = 8'b00000000;	//         
        11'he359: data = 8'b00000000;	//         
        11'he35a: data = 8'b00000000;	//         
        11'he35b: data = 8'b00000000;	//         
        11'he35c: data = 8'b00000000;	//         
        11'he35d: data = 8'b00000000;	//         
        11'he35e: data = 8'b00000000;	//         
        11'he35f: data = 8'b00000000;	//         

    // code xe36 (ึ)
        11'he360: data = 8'b00000000;	//         
        11'he361: data = 8'b00000000;	//         
        11'he362: data = 8'b00000000;	//         
        11'he363: data = 8'b00000011;	//       **
        11'he364: data = 8'b00001111;	//     ****
        11'he365: data = 8'b00000000;	//         
        11'he366: data = 8'b00000000;	//         
        11'he367: data = 8'b00000000;	//         
        11'he368: data = 8'b00000000;	//         
        11'he369: data = 8'b00000000;	//         
        11'he36a: data = 8'b00000000;	//         
        11'he36b: data = 8'b00000000;	//         
        11'he36c: data = 8'b00000000;	//         
        11'he36d: data = 8'b00000000;	//         
        11'he36e: data = 8'b00000000;	//         
        11'he36f: data = 8'b00000000;	//         

    // code xe37 (ื)
        11'he370: data = 8'b00000000;	//         
        11'he371: data = 8'b00000000;	//         
        11'he372: data = 8'b00000000;	//         
        11'he373: data = 8'b00000000;	//         
        11'he374: data = 8'b00001111;	//     ****
        11'he375: data = 8'b00000000;	//         
        11'he376: data = 8'b00000000;	//         
        11'he377: data = 8'b00000000;	//         
        11'he378: data = 8'b00000000;	//         
        11'he379: data = 8'b00000000;	//         
        11'he37a: data = 8'b00000000;	//         
        11'he37b: data = 8'b00000000;	//         
        11'he37c: data = 8'b00000000;	//         
        11'he37d: data = 8'b00000000;	//         
        11'he37e: data = 8'b00000000;	//         
        11'he37f: data = 8'b00000000;	//         

    // code xe38 (ุ)
        11'he380: data = 8'b00000000;	//         
        11'he381: data = 8'b00000000;	//         
        11'he382: data = 8'b00000000;	//         
        11'he383: data = 8'b00000000;	//         
        11'he384: data = 8'b00000000;	//         
        11'he385: data = 8'b00000000;	//         
        11'he386: data = 8'b00000000;	//         
        11'he387: data = 8'b00000000;	//         
        11'he388: data = 8'b00000000;	//         
        11'he389: data = 8'b00000000;	//         
        11'he38a: data = 8'b00000000;	//         
        11'he38b: data = 8'b00000001;	//        *
        11'he38c: data = 8'b00000001;	//        *
        11'he38d: data = 8'b00000000;	//         
        11'he38e: data = 8'b00000000;	//         
        11'he38f: data = 8'b00000000;	//         

    // code xe39 (ู)
        11'he390: data = 8'b00000000;	//         
        11'he391: data = 8'b00000000;	//         
        11'he392: data = 8'b00000000;	//         
        11'he393: data = 8'b00000000;	//         
        11'he394: data = 8'b00000000;	//         
        11'he395: data = 8'b00000000;	//         
        11'he396: data = 8'b00000000;	//         
        11'he397: data = 8'b00000000;	//         
        11'he398: data = 8'b00000000;	//         
        11'he399: data = 8'b00000000;	//         
        11'he39a: data = 8'b00000000;	//         
        11'he39b: data = 8'b00001001;	//     *  *
        11'he39c: data = 8'b00001111;	//     ****
        11'he39d: data = 8'b00000000;	//         
        11'he39e: data = 8'b00000000;	//         
        11'he39f: data = 8'b00000000;	//         

    // code xe40 (เ)
        11'he400: data = 8'b00000000;	//         
        11'he401: data = 8'b00000000;	//         
        11'he402: data = 8'b00000000;	//         
        11'he403: data = 8'b11000000;	// **      
        11'he404: data = 8'b11000000;	// **      
        11'he405: data = 8'b11000000;	// **      
        11'he406: data = 8'b11000000;	// **      
        11'he407: data = 8'b11000000;	// **      
        11'he408: data = 8'b11000000;	// **      
        11'he409: data = 8'b11000000;	// **      
        11'he40a: data = 8'b00000000;	//         
        11'he40b: data = 8'b00000000;	//         
        11'he40c: data = 8'b00000000;	//         
        11'he40d: data = 8'b00000000;	//         
        11'he40e: data = 8'b00000000;	//         
        11'he40f: data = 8'b00000000;	//         

    // code xe41 (แ)
        11'he410: data = 8'b00000000;	//         
        11'he411: data = 8'b00000000;	//         
        11'he412: data = 8'b00000000;	//         
        11'he413: data = 8'b11001000;	// **  *   
        11'he414: data = 8'b11001000;	// **  *   
        11'he415: data = 8'b11001000;	// **  *   
        11'he416: data = 8'b11001000;	// **  *   
        11'he417: data = 8'b11001000;	// **  *   
        11'he418: data = 8'b11001000;	// **  *   
        11'he419: data = 8'b11001000;	// **  *   
        11'he41a: data = 8'b00000000;	//         
        11'he41b: data = 8'b00000000;	//         
        11'he41c: data = 8'b00000000;	//         
        11'he41d: data = 8'b00000000;	//         
        11'he41e: data = 8'b00000000;	//         
        11'he41f: data = 8'b00000000;	//         

    // code xe42 (โ)
        11'he420: data = 8'b10000000;	// *       
        11'he421: data = 8'b11000000;	// **      
        11'he422: data = 8'b11000000;	// **      
        11'he423: data = 8'b11000000;	// **      
        11'he424: data = 8'b11000000;	// **      
        11'he425: data = 8'b11000000;	// **      
        11'he426: data = 8'b11000000;	// **      
        11'he427: data = 8'b11000000;	// **      
        11'he428: data = 8'b11000000;	// **      
        11'he429: data = 8'b11000000;	// **      
        11'he42a: data = 8'b00000000;	//         
        11'he42b: data = 8'b00000000;	//         
        11'he42c: data = 8'b00000000;	//         
        11'he42d: data = 8'b00000000;	//         
        11'he42e: data = 8'b00000000;	//         
        11'he42f: data = 8'b00000000;	//         

    // code xe43 (ใ)
        11'he430: data = 8'b11000000;	// **      
        11'he431: data = 8'b11000000;	// **      
        11'he432: data = 8'b11000000;	// **      
        11'he433: data = 8'b11000000;	// **      
        11'he434: data = 8'b11000000;	// **      
        11'he435: data = 8'b11000000;	// **      
        11'he436: data = 8'b11000000;	// **      
        11'he437: data = 8'b11000000;	// **      
        11'he438: data = 8'b11000000;	// **      
        11'he439: data = 8'b11000000;	// **      
        11'he43a: data = 8'b00000000;	//         
        11'he43b: data = 8'b00000000;	//         
        11'he43c: data = 8'b00000000;	//         
        11'he43d: data = 8'b00000000;	//         
        11'he43e: data = 8'b00000000;	//         
        11'he43f: data = 8'b00000000;	//         

    // code xe44 (ไ)
        11'he440: data = 8'b11000000;	// **      
        11'he441: data = 8'b11000000;	// **      
        11'he442: data = 8'b11000000;	// **      
        11'he443: data = 8'b11000000;	// **      
        11'he444: data = 8'b11000000;	// **      
        11'he445: data = 8'b11000000;	// **      
        11'he446: data = 8'b11000000;	// **      
        11'he447: data = 8'b11000000;	// **      
        11'he448: data = 8'b11000000;	// **      
        11'he449: data = 8'b11000000;	// **      
        11'he44a: data = 8'b00000000;	//         
        11'he44b: data = 8'b00000000;	//         
        11'he44c: data = 8'b00000000;	//         
        11'he44d: data = 8'b00000000;	//         
        11'he44e: data = 8'b00000000;	//         
        11'he44f: data = 8'b00000000;	//         

            default: data = 8'b00000000; // Default to zero
        endcase
 endmodule
    